library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity sincos_lut is
generic(
  N : integer := 16
);
port
(
  reset           : in  std_logic;
  clk             : in  std_logic;
  clk_en          : in  std_logic;
  theta           : in  std_logic_vector(11 downto 0);
  sin_data        : out std_logic_vector(N-1 downto 0);
  cos_data        : out std_logic_vector(N-1 downto 0)
);
end sincos_lut;

architecture rtl of sincos_lut is

  signal theta_int      : integer range 0 to 4095 := 0;
  signal sin_data_int   : unsigned(N-1 downto 0);
  signal cos_data_int   : unsigned(N-1 downto 0);

  signal negate : std_logic := '0';

begin

  process(clk)
  begin
    if rising_edge(clk) then
      if (to_integer(unsigned(theta)) > 2047) then
        theta_int <= 4095 - to_integer(unsigned(theta));
        negate <= '1';
      else
        theta_int <= to_integer(unsigned(theta));
        negate <= '0';
      end if;
    end if;
  end process;

  process(reset,clk)
  begin
    if(reset = '1')then
      sin_data_int <= to_unsigned(0,N);
      cos_data_int <= to_unsigned(0,N);
    elsif(rising_edge(clk)) then
      if clk_en = '1' then
        if (negate = '1') then
          sin_data <= std_logic_vector(not(sin_data_int) + 1);
          cos_data <= std_logic_vector(cos_data_int);
        else
          sin_data <= std_logic_vector(sin_data_int);
          cos_data <= std_logic_vector(cos_data_int);
        end if;

        case theta_int is
          when 0 =>   sin_data_int <= to_unsigned(0,N); cos_data_int <= to_unsigned(16384,N);
          when 1 =>   sin_data_int <= to_unsigned(25,N); cos_data_int <= to_unsigned(16383,N);
          when 2 =>   sin_data_int <= to_unsigned(50,N); cos_data_int <= to_unsigned(16383,N);
          when 3 =>   sin_data_int <= to_unsigned(75,N); cos_data_int <= to_unsigned(16383,N);
          when 4 =>   sin_data_int <= to_unsigned(100,N); cos_data_int <= to_unsigned(16383,N);
          when 5 =>   sin_data_int <= to_unsigned(125,N); cos_data_int <= to_unsigned(16383,N);
          when 6 =>   sin_data_int <= to_unsigned(150,N); cos_data_int <= to_unsigned(16383,N);
          when 7 =>   sin_data_int <= to_unsigned(175,N); cos_data_int <= to_unsigned(16383,N);
          when 8 =>   sin_data_int <= to_unsigned(201,N); cos_data_int <= to_unsigned(16382,N);
          when 9 =>   sin_data_int <= to_unsigned(226,N); cos_data_int <= to_unsigned(16382,N);
          when 10 =>   sin_data_int <= to_unsigned(251,N); cos_data_int <= to_unsigned(16382,N);
          when 11 =>   sin_data_int <= to_unsigned(276,N); cos_data_int <= to_unsigned(16381,N);
          when 12 =>   sin_data_int <= to_unsigned(301,N); cos_data_int <= to_unsigned(16381,N);
          when 13 =>   sin_data_int <= to_unsigned(326,N); cos_data_int <= to_unsigned(16380,N);
          when 14 =>   sin_data_int <= to_unsigned(351,N); cos_data_int <= to_unsigned(16380,N);
          when 15 =>   sin_data_int <= to_unsigned(376,N); cos_data_int <= to_unsigned(16379,N);
          when 16 =>   sin_data_int <= to_unsigned(402,N); cos_data_int <= to_unsigned(16379,N);
          when 17 =>   sin_data_int <= to_unsigned(427,N); cos_data_int <= to_unsigned(16378,N);
          when 18 =>   sin_data_int <= to_unsigned(452,N); cos_data_int <= to_unsigned(16377,N);
          when 19 =>   sin_data_int <= to_unsigned(477,N); cos_data_int <= to_unsigned(16377,N);
          when 20 =>   sin_data_int <= to_unsigned(502,N); cos_data_int <= to_unsigned(16376,N);
          when 21 =>   sin_data_int <= to_unsigned(527,N); cos_data_int <= to_unsigned(16375,N);
          when 22 =>   sin_data_int <= to_unsigned(552,N); cos_data_int <= to_unsigned(16374,N);
          when 23 =>   sin_data_int <= to_unsigned(577,N); cos_data_int <= to_unsigned(16373,N);
          when 24 =>   sin_data_int <= to_unsigned(603,N); cos_data_int <= to_unsigned(16372,N);
          when 25 =>   sin_data_int <= to_unsigned(628,N); cos_data_int <= to_unsigned(16371,N);
          when 26 =>   sin_data_int <= to_unsigned(653,N); cos_data_int <= to_unsigned(16370,N);
          when 27 =>   sin_data_int <= to_unsigned(678,N); cos_data_int <= to_unsigned(16369,N);
          when 28 =>   sin_data_int <= to_unsigned(703,N); cos_data_int <= to_unsigned(16368,N);
          when 29 =>   sin_data_int <= to_unsigned(728,N); cos_data_int <= to_unsigned(16367,N);
          when 30 =>   sin_data_int <= to_unsigned(753,N); cos_data_int <= to_unsigned(16366,N);
          when 31 =>   sin_data_int <= to_unsigned(778,N); cos_data_int <= to_unsigned(16365,N);
          when 32 =>   sin_data_int <= to_unsigned(803,N); cos_data_int <= to_unsigned(16364,N);
          when 33 =>   sin_data_int <= to_unsigned(829,N); cos_data_int <= to_unsigned(16363,N);
          when 34 =>   sin_data_int <= to_unsigned(854,N); cos_data_int <= to_unsigned(16361,N);
          when 35 =>   sin_data_int <= to_unsigned(879,N); cos_data_int <= to_unsigned(16360,N);
          when 36 =>   sin_data_int <= to_unsigned(904,N); cos_data_int <= to_unsigned(16359,N);
          when 37 =>   sin_data_int <= to_unsigned(929,N); cos_data_int <= to_unsigned(16357,N);
          when 38 =>   sin_data_int <= to_unsigned(954,N); cos_data_int <= to_unsigned(16356,N);
          when 39 =>   sin_data_int <= to_unsigned(979,N); cos_data_int <= to_unsigned(16354,N);
          when 40 =>   sin_data_int <= to_unsigned(1004,N); cos_data_int <= to_unsigned(16353,N);
          when 41 =>   sin_data_int <= to_unsigned(1029,N); cos_data_int <= to_unsigned(16351,N);
          when 42 =>   sin_data_int <= to_unsigned(1054,N); cos_data_int <= to_unsigned(16350,N);
          when 43 =>   sin_data_int <= to_unsigned(1079,N); cos_data_int <= to_unsigned(16348,N);
          when 44 =>   sin_data_int <= to_unsigned(1105,N); cos_data_int <= to_unsigned(16346,N);
          when 45 =>   sin_data_int <= to_unsigned(1130,N); cos_data_int <= to_unsigned(16344,N);
          when 46 =>   sin_data_int <= to_unsigned(1155,N); cos_data_int <= to_unsigned(16343,N);
          when 47 =>   sin_data_int <= to_unsigned(1180,N); cos_data_int <= to_unsigned(16341,N);
          when 48 =>   sin_data_int <= to_unsigned(1205,N); cos_data_int <= to_unsigned(16339,N);
          when 49 =>   sin_data_int <= to_unsigned(1230,N); cos_data_int <= to_unsigned(16337,N);
          when 50 =>   sin_data_int <= to_unsigned(1255,N); cos_data_int <= to_unsigned(16335,N);
          when 51 =>   sin_data_int <= to_unsigned(1280,N); cos_data_int <= to_unsigned(16333,N);
          when 52 =>   sin_data_int <= to_unsigned(1305,N); cos_data_int <= to_unsigned(16331,N);
          when 53 =>   sin_data_int <= to_unsigned(1330,N); cos_data_int <= to_unsigned(16329,N);
          when 54 =>   sin_data_int <= to_unsigned(1355,N); cos_data_int <= to_unsigned(16327,N);
          when 55 =>   sin_data_int <= to_unsigned(1380,N); cos_data_int <= to_unsigned(16325,N);
          when 56 =>   sin_data_int <= to_unsigned(1405,N); cos_data_int <= to_unsigned(16323,N);
          when 57 =>   sin_data_int <= to_unsigned(1430,N); cos_data_int <= to_unsigned(16321,N);
          when 58 =>   sin_data_int <= to_unsigned(1455,N); cos_data_int <= to_unsigned(16319,N);
          when 59 =>   sin_data_int <= to_unsigned(1480,N); cos_data_int <= to_unsigned(16316,N);
          when 60 =>   sin_data_int <= to_unsigned(1505,N); cos_data_int <= to_unsigned(16314,N);
          when 61 =>   sin_data_int <= to_unsigned(1530,N); cos_data_int <= to_unsigned(16312,N);
          when 62 =>   sin_data_int <= to_unsigned(1555,N); cos_data_int <= to_unsigned(16309,N);
          when 63 =>   sin_data_int <= to_unsigned(1580,N); cos_data_int <= to_unsigned(16307,N);
          when 64 =>   sin_data_int <= to_unsigned(1605,N); cos_data_int <= to_unsigned(16305,N);
          when 65 =>   sin_data_int <= to_unsigned(1630,N); cos_data_int <= to_unsigned(16302,N);
          when 66 =>   sin_data_int <= to_unsigned(1655,N); cos_data_int <= to_unsigned(16300,N);
          when 67 =>   sin_data_int <= to_unsigned(1680,N); cos_data_int <= to_unsigned(16297,N);
          when 68 =>   sin_data_int <= to_unsigned(1705,N); cos_data_int <= to_unsigned(16294,N);
          when 69 =>   sin_data_int <= to_unsigned(1730,N); cos_data_int <= to_unsigned(16292,N);
          when 70 =>   sin_data_int <= to_unsigned(1755,N); cos_data_int <= to_unsigned(16289,N);
          when 71 =>   sin_data_int <= to_unsigned(1780,N); cos_data_int <= to_unsigned(16286,N);
          when 72 =>   sin_data_int <= to_unsigned(1805,N); cos_data_int <= to_unsigned(16284,N);
          when 73 =>   sin_data_int <= to_unsigned(1830,N); cos_data_int <= to_unsigned(16281,N);
          when 74 =>   sin_data_int <= to_unsigned(1855,N); cos_data_int <= to_unsigned(16278,N);
          when 75 =>   sin_data_int <= to_unsigned(1880,N); cos_data_int <= to_unsigned(16275,N);
          when 76 =>   sin_data_int <= to_unsigned(1905,N); cos_data_int <= to_unsigned(16272,N);
          when 77 =>   sin_data_int <= to_unsigned(1930,N); cos_data_int <= to_unsigned(16269,N);
          when 78 =>   sin_data_int <= to_unsigned(1955,N); cos_data_int <= to_unsigned(16266,N);
          when 79 =>   sin_data_int <= to_unsigned(1980,N); cos_data_int <= to_unsigned(16263,N);
          when 80 =>   sin_data_int <= to_unsigned(2005,N); cos_data_int <= to_unsigned(16260,N);
          when 81 =>   sin_data_int <= to_unsigned(2030,N); cos_data_int <= to_unsigned(16257,N);
          when 82 =>   sin_data_int <= to_unsigned(2055,N); cos_data_int <= to_unsigned(16254,N);
          when 83 =>   sin_data_int <= to_unsigned(2080,N); cos_data_int <= to_unsigned(16251,N);
          when 84 =>   sin_data_int <= to_unsigned(2105,N); cos_data_int <= to_unsigned(16248,N);
          when 85 =>   sin_data_int <= to_unsigned(2130,N); cos_data_int <= to_unsigned(16244,N);
          when 86 =>   sin_data_int <= to_unsigned(2155,N); cos_data_int <= to_unsigned(16241,N);
          when 87 =>   sin_data_int <= to_unsigned(2180,N); cos_data_int <= to_unsigned(16238,N);
          when 88 =>   sin_data_int <= to_unsigned(2204,N); cos_data_int <= to_unsigned(16234,N);
          when 89 =>   sin_data_int <= to_unsigned(2229,N); cos_data_int <= to_unsigned(16231,N);
          when 90 =>   sin_data_int <= to_unsigned(2254,N); cos_data_int <= to_unsigned(16228,N);
          when 91 =>   sin_data_int <= to_unsigned(2279,N); cos_data_int <= to_unsigned(16224,N);
          when 92 =>   sin_data_int <= to_unsigned(2304,N); cos_data_int <= to_unsigned(16221,N);
          when 93 =>   sin_data_int <= to_unsigned(2329,N); cos_data_int <= to_unsigned(16217,N);
          when 94 =>   sin_data_int <= to_unsigned(2354,N); cos_data_int <= to_unsigned(16213,N);
          when 95 =>   sin_data_int <= to_unsigned(2379,N); cos_data_int <= to_unsigned(16210,N);
          when 96 =>   sin_data_int <= to_unsigned(2404,N); cos_data_int <= to_unsigned(16206,N);
          when 97 =>   sin_data_int <= to_unsigned(2428,N); cos_data_int <= to_unsigned(16202,N);
          when 98 =>   sin_data_int <= to_unsigned(2453,N); cos_data_int <= to_unsigned(16199,N);
          when 99 =>   sin_data_int <= to_unsigned(2478,N); cos_data_int <= to_unsigned(16195,N);
          when 100 =>   sin_data_int <= to_unsigned(2503,N); cos_data_int <= to_unsigned(16191,N);
          when 101 =>   sin_data_int <= to_unsigned(2528,N); cos_data_int <= to_unsigned(16187,N);
          when 102 =>   sin_data_int <= to_unsigned(2553,N); cos_data_int <= to_unsigned(16183,N);
          when 103 =>   sin_data_int <= to_unsigned(2577,N); cos_data_int <= to_unsigned(16179,N);
          when 104 =>   sin_data_int <= to_unsigned(2602,N); cos_data_int <= to_unsigned(16175,N);
          when 105 =>   sin_data_int <= to_unsigned(2627,N); cos_data_int <= to_unsigned(16171,N);
          when 106 =>   sin_data_int <= to_unsigned(2652,N); cos_data_int <= to_unsigned(16167,N);
          when 107 =>   sin_data_int <= to_unsigned(2677,N); cos_data_int <= to_unsigned(16163,N);
          when 108 =>   sin_data_int <= to_unsigned(2701,N); cos_data_int <= to_unsigned(16159,N);
          when 109 =>   sin_data_int <= to_unsigned(2726,N); cos_data_int <= to_unsigned(16155,N);
          when 110 =>   sin_data_int <= to_unsigned(2751,N); cos_data_int <= to_unsigned(16151,N);
          when 111 =>   sin_data_int <= to_unsigned(2776,N); cos_data_int <= to_unsigned(16147,N);
          when 112 =>   sin_data_int <= to_unsigned(2801,N); cos_data_int <= to_unsigned(16142,N);
          when 113 =>   sin_data_int <= to_unsigned(2825,N); cos_data_int <= to_unsigned(16138,N);
          when 114 =>   sin_data_int <= to_unsigned(2850,N); cos_data_int <= to_unsigned(16134,N);
          when 115 =>   sin_data_int <= to_unsigned(2875,N); cos_data_int <= to_unsigned(16129,N);
          when 116 =>   sin_data_int <= to_unsigned(2900,N); cos_data_int <= to_unsigned(16125,N);
          when 117 =>   sin_data_int <= to_unsigned(2924,N); cos_data_int <= to_unsigned(16120,N);
          when 118 =>   sin_data_int <= to_unsigned(2949,N); cos_data_int <= to_unsigned(16116,N);
          when 119 =>   sin_data_int <= to_unsigned(2974,N); cos_data_int <= to_unsigned(16111,N);
          when 120 =>   sin_data_int <= to_unsigned(2998,N); cos_data_int <= to_unsigned(16107,N);
          when 121 =>   sin_data_int <= to_unsigned(3023,N); cos_data_int <= to_unsigned(16102,N);
          when 122 =>   sin_data_int <= to_unsigned(3048,N); cos_data_int <= to_unsigned(16097,N);
          when 123 =>   sin_data_int <= to_unsigned(3073,N); cos_data_int <= to_unsigned(16093,N);
          when 124 =>   sin_data_int <= to_unsigned(3097,N); cos_data_int <= to_unsigned(16088,N);
          when 125 =>   sin_data_int <= to_unsigned(3122,N); cos_data_int <= to_unsigned(16083,N);
          when 126 =>   sin_data_int <= to_unsigned(3147,N); cos_data_int <= to_unsigned(16078,N);
          when 127 =>   sin_data_int <= to_unsigned(3171,N); cos_data_int <= to_unsigned(16074,N);
          when 128 =>   sin_data_int <= to_unsigned(3196,N); cos_data_int <= to_unsigned(16069,N);
          when 129 =>   sin_data_int <= to_unsigned(3221,N); cos_data_int <= to_unsigned(16064,N);
          when 130 =>   sin_data_int <= to_unsigned(3245,N); cos_data_int <= to_unsigned(16059,N);
          when 131 =>   sin_data_int <= to_unsigned(3270,N); cos_data_int <= to_unsigned(16054,N);
          when 132 =>   sin_data_int <= to_unsigned(3294,N); cos_data_int <= to_unsigned(16049,N);
          when 133 =>   sin_data_int <= to_unsigned(3319,N); cos_data_int <= to_unsigned(16044,N);
          when 134 =>   sin_data_int <= to_unsigned(3344,N); cos_data_int <= to_unsigned(16039,N);
          when 135 =>   sin_data_int <= to_unsigned(3368,N); cos_data_int <= to_unsigned(16033,N);
          when 136 =>   sin_data_int <= to_unsigned(3393,N); cos_data_int <= to_unsigned(16028,N);
          when 137 =>   sin_data_int <= to_unsigned(3417,N); cos_data_int <= to_unsigned(16023,N);
          when 138 =>   sin_data_int <= to_unsigned(3442,N); cos_data_int <= to_unsigned(16018,N);
          when 139 =>   sin_data_int <= to_unsigned(3467,N); cos_data_int <= to_unsigned(16012,N);
          when 140 =>   sin_data_int <= to_unsigned(3491,N); cos_data_int <= to_unsigned(16007,N);
          when 141 =>   sin_data_int <= to_unsigned(3516,N); cos_data_int <= to_unsigned(16002,N);
          when 142 =>   sin_data_int <= to_unsigned(3540,N); cos_data_int <= to_unsigned(15996,N);
          when 143 =>   sin_data_int <= to_unsigned(3565,N); cos_data_int <= to_unsigned(15991,N);
          when 144 =>   sin_data_int <= to_unsigned(3589,N); cos_data_int <= to_unsigned(15985,N);
          when 145 =>   sin_data_int <= to_unsigned(3614,N); cos_data_int <= to_unsigned(15980,N);
          when 146 =>   sin_data_int <= to_unsigned(3638,N); cos_data_int <= to_unsigned(15974,N);
          when 147 =>   sin_data_int <= to_unsigned(3663,N); cos_data_int <= to_unsigned(15969,N);
          when 148 =>   sin_data_int <= to_unsigned(3687,N); cos_data_int <= to_unsigned(15963,N);
          when 149 =>   sin_data_int <= to_unsigned(3712,N); cos_data_int <= to_unsigned(15957,N);
          when 150 =>   sin_data_int <= to_unsigned(3736,N); cos_data_int <= to_unsigned(15952,N);
          when 151 =>   sin_data_int <= to_unsigned(3761,N); cos_data_int <= to_unsigned(15946,N);
          when 152 =>   sin_data_int <= to_unsigned(3785,N); cos_data_int <= to_unsigned(15940,N);
          when 153 =>   sin_data_int <= to_unsigned(3810,N); cos_data_int <= to_unsigned(15934,N);
          when 154 =>   sin_data_int <= to_unsigned(3834,N); cos_data_int <= to_unsigned(15928,N);
          when 155 =>   sin_data_int <= to_unsigned(3858,N); cos_data_int <= to_unsigned(15923,N);
          when 156 =>   sin_data_int <= to_unsigned(3883,N); cos_data_int <= to_unsigned(15917,N);
          when 157 =>   sin_data_int <= to_unsigned(3907,N); cos_data_int <= to_unsigned(15911,N);
          when 158 =>   sin_data_int <= to_unsigned(3932,N); cos_data_int <= to_unsigned(15905,N);
          when 159 =>   sin_data_int <= to_unsigned(3956,N); cos_data_int <= to_unsigned(15899,N);
          when 160 =>   sin_data_int <= to_unsigned(3980,N); cos_data_int <= to_unsigned(15892,N);
          when 161 =>   sin_data_int <= to_unsigned(4005,N); cos_data_int <= to_unsigned(15886,N);
          when 162 =>   sin_data_int <= to_unsigned(4029,N); cos_data_int <= to_unsigned(15880,N);
          when 163 =>   sin_data_int <= to_unsigned(4054,N); cos_data_int <= to_unsigned(15874,N);
          when 164 =>   sin_data_int <= to_unsigned(4078,N); cos_data_int <= to_unsigned(15868,N);
          when 165 =>   sin_data_int <= to_unsigned(4102,N); cos_data_int <= to_unsigned(15861,N);
          when 166 =>   sin_data_int <= to_unsigned(4127,N); cos_data_int <= to_unsigned(15855,N);
          when 167 =>   sin_data_int <= to_unsigned(4151,N); cos_data_int <= to_unsigned(15849,N);
          when 168 =>   sin_data_int <= to_unsigned(4175,N); cos_data_int <= to_unsigned(15842,N);
          when 169 =>   sin_data_int <= to_unsigned(4200,N); cos_data_int <= to_unsigned(15836,N);
          when 170 =>   sin_data_int <= to_unsigned(4224,N); cos_data_int <= to_unsigned(15830,N);
          when 171 =>   sin_data_int <= to_unsigned(4248,N); cos_data_int <= to_unsigned(15823,N);
          when 172 =>   sin_data_int <= to_unsigned(4272,N); cos_data_int <= to_unsigned(15817,N);
          when 173 =>   sin_data_int <= to_unsigned(4297,N); cos_data_int <= to_unsigned(15810,N);
          when 174 =>   sin_data_int <= to_unsigned(4321,N); cos_data_int <= to_unsigned(15803,N);
          when 175 =>   sin_data_int <= to_unsigned(4345,N); cos_data_int <= to_unsigned(15797,N);
          when 176 =>   sin_data_int <= to_unsigned(4369,N); cos_data_int <= to_unsigned(15790,N);
          when 177 =>   sin_data_int <= to_unsigned(4394,N); cos_data_int <= to_unsigned(15783,N);
          when 178 =>   sin_data_int <= to_unsigned(4418,N); cos_data_int <= to_unsigned(15777,N);
          when 179 =>   sin_data_int <= to_unsigned(4442,N); cos_data_int <= to_unsigned(15770,N);
          when 180 =>   sin_data_int <= to_unsigned(4466,N); cos_data_int <= to_unsigned(15763,N);
          when 181 =>   sin_data_int <= to_unsigned(4490,N); cos_data_int <= to_unsigned(15756,N);
          when 182 =>   sin_data_int <= to_unsigned(4514,N); cos_data_int <= to_unsigned(15749,N);
          when 183 =>   sin_data_int <= to_unsigned(4539,N); cos_data_int <= to_unsigned(15742,N);
          when 184 =>   sin_data_int <= to_unsigned(4563,N); cos_data_int <= to_unsigned(15735,N);
          when 185 =>   sin_data_int <= to_unsigned(4587,N); cos_data_int <= to_unsigned(15728,N);
          when 186 =>   sin_data_int <= to_unsigned(4611,N); cos_data_int <= to_unsigned(15721,N);
          when 187 =>   sin_data_int <= to_unsigned(4635,N); cos_data_int <= to_unsigned(15714,N);
          when 188 =>   sin_data_int <= to_unsigned(4659,N); cos_data_int <= to_unsigned(15707,N);
          when 189 =>   sin_data_int <= to_unsigned(4683,N); cos_data_int <= to_unsigned(15700,N);
          when 190 =>   sin_data_int <= to_unsigned(4707,N); cos_data_int <= to_unsigned(15693,N);
          when 191 =>   sin_data_int <= to_unsigned(4731,N); cos_data_int <= to_unsigned(15685,N);
          when 192 =>   sin_data_int <= to_unsigned(4756,N); cos_data_int <= to_unsigned(15678,N);
          when 193 =>   sin_data_int <= to_unsigned(4780,N); cos_data_int <= to_unsigned(15671,N);
          when 194 =>   sin_data_int <= to_unsigned(4804,N); cos_data_int <= to_unsigned(15663,N);
          when 195 =>   sin_data_int <= to_unsigned(4828,N); cos_data_int <= to_unsigned(15656,N);
          when 196 =>   sin_data_int <= to_unsigned(4852,N); cos_data_int <= to_unsigned(15649,N);
          when 197 =>   sin_data_int <= to_unsigned(4876,N); cos_data_int <= to_unsigned(15641,N);
          when 198 =>   sin_data_int <= to_unsigned(4900,N); cos_data_int <= to_unsigned(15634,N);
          when 199 =>   sin_data_int <= to_unsigned(4924,N); cos_data_int <= to_unsigned(15626,N);
          when 200 =>   sin_data_int <= to_unsigned(4948,N); cos_data_int <= to_unsigned(15618,N);
          when 201 =>   sin_data_int <= to_unsigned(4972,N); cos_data_int <= to_unsigned(15611,N);
          when 202 =>   sin_data_int <= to_unsigned(4995,N); cos_data_int <= to_unsigned(15603,N);
          when 203 =>   sin_data_int <= to_unsigned(5019,N); cos_data_int <= to_unsigned(15596,N);
          when 204 =>   sin_data_int <= to_unsigned(5043,N); cos_data_int <= to_unsigned(15588,N);
          when 205 =>   sin_data_int <= to_unsigned(5067,N); cos_data_int <= to_unsigned(15580,N);
          when 206 =>   sin_data_int <= to_unsigned(5091,N); cos_data_int <= to_unsigned(15572,N);
          when 207 =>   sin_data_int <= to_unsigned(5115,N); cos_data_int <= to_unsigned(15564,N);
          when 208 =>   sin_data_int <= to_unsigned(5139,N); cos_data_int <= to_unsigned(15557,N);
          when 209 =>   sin_data_int <= to_unsigned(5163,N); cos_data_int <= to_unsigned(15549,N);
          when 210 =>   sin_data_int <= to_unsigned(5187,N); cos_data_int <= to_unsigned(15541,N);
          when 211 =>   sin_data_int <= to_unsigned(5210,N); cos_data_int <= to_unsigned(15533,N);
          when 212 =>   sin_data_int <= to_unsigned(5234,N); cos_data_int <= to_unsigned(15525,N);
          when 213 =>   sin_data_int <= to_unsigned(5258,N); cos_data_int <= to_unsigned(15517,N);
          when 214 =>   sin_data_int <= to_unsigned(5282,N); cos_data_int <= to_unsigned(15509,N);
          when 215 =>   sin_data_int <= to_unsigned(5306,N); cos_data_int <= to_unsigned(15500,N);
          when 216 =>   sin_data_int <= to_unsigned(5329,N); cos_data_int <= to_unsigned(15492,N);
          when 217 =>   sin_data_int <= to_unsigned(5353,N); cos_data_int <= to_unsigned(15484,N);
          when 218 =>   sin_data_int <= to_unsigned(5377,N); cos_data_int <= to_unsigned(15476,N);
          when 219 =>   sin_data_int <= to_unsigned(5401,N); cos_data_int <= to_unsigned(15468,N);
          when 220 =>   sin_data_int <= to_unsigned(5424,N); cos_data_int <= to_unsigned(15459,N);
          when 221 =>   sin_data_int <= to_unsigned(5448,N); cos_data_int <= to_unsigned(15451,N);
          when 222 =>   sin_data_int <= to_unsigned(5472,N); cos_data_int <= to_unsigned(15443,N);
          when 223 =>   sin_data_int <= to_unsigned(5495,N); cos_data_int <= to_unsigned(15434,N);
          when 224 =>   sin_data_int <= to_unsigned(5519,N); cos_data_int <= to_unsigned(15426,N);
          when 225 =>   sin_data_int <= to_unsigned(5543,N); cos_data_int <= to_unsigned(15417,N);
          when 226 =>   sin_data_int <= to_unsigned(5566,N); cos_data_int <= to_unsigned(15409,N);
          when 227 =>   sin_data_int <= to_unsigned(5590,N); cos_data_int <= to_unsigned(15400,N);
          when 228 =>   sin_data_int <= to_unsigned(5614,N); cos_data_int <= to_unsigned(15392,N);
          when 229 =>   sin_data_int <= to_unsigned(5637,N); cos_data_int <= to_unsigned(15383,N);
          when 230 =>   sin_data_int <= to_unsigned(5661,N); cos_data_int <= to_unsigned(15374,N);
          when 231 =>   sin_data_int <= to_unsigned(5684,N); cos_data_int <= to_unsigned(15366,N);
          when 232 =>   sin_data_int <= to_unsigned(5708,N); cos_data_int <= to_unsigned(15357,N);
          when 233 =>   sin_data_int <= to_unsigned(5732,N); cos_data_int <= to_unsigned(15348,N);
          when 234 =>   sin_data_int <= to_unsigned(5755,N); cos_data_int <= to_unsigned(15339,N);
          when 235 =>   sin_data_int <= to_unsigned(5779,N); cos_data_int <= to_unsigned(15330,N);
          when 236 =>   sin_data_int <= to_unsigned(5802,N); cos_data_int <= to_unsigned(15322,N);
          when 237 =>   sin_data_int <= to_unsigned(5826,N); cos_data_int <= to_unsigned(15313,N);
          when 238 =>   sin_data_int <= to_unsigned(5849,N); cos_data_int <= to_unsigned(15304,N);
          when 239 =>   sin_data_int <= to_unsigned(5873,N); cos_data_int <= to_unsigned(15295,N);
          when 240 =>   sin_data_int <= to_unsigned(5896,N); cos_data_int <= to_unsigned(15286,N);
          when 241 =>   sin_data_int <= to_unsigned(5919,N); cos_data_int <= to_unsigned(15277,N);
          when 242 =>   sin_data_int <= to_unsigned(5943,N); cos_data_int <= to_unsigned(15267,N);
          when 243 =>   sin_data_int <= to_unsigned(5966,N); cos_data_int <= to_unsigned(15258,N);
          when 244 =>   sin_data_int <= to_unsigned(5990,N); cos_data_int <= to_unsigned(15249,N);
          when 245 =>   sin_data_int <= to_unsigned(6013,N); cos_data_int <= to_unsigned(15240,N);
          when 246 =>   sin_data_int <= to_unsigned(6036,N); cos_data_int <= to_unsigned(15231,N);
          when 247 =>   sin_data_int <= to_unsigned(6060,N); cos_data_int <= to_unsigned(15221,N);
          when 248 =>   sin_data_int <= to_unsigned(6083,N); cos_data_int <= to_unsigned(15212,N);
          when 249 =>   sin_data_int <= to_unsigned(6106,N); cos_data_int <= to_unsigned(15203,N);
          when 250 =>   sin_data_int <= to_unsigned(6130,N); cos_data_int <= to_unsigned(15193,N);
          when 251 =>   sin_data_int <= to_unsigned(6153,N); cos_data_int <= to_unsigned(15184,N);
          when 252 =>   sin_data_int <= to_unsigned(6176,N); cos_data_int <= to_unsigned(15175,N);
          when 253 =>   sin_data_int <= to_unsigned(6200,N); cos_data_int <= to_unsigned(15165,N);
          when 254 =>   sin_data_int <= to_unsigned(6223,N); cos_data_int <= to_unsigned(15156,N);
          when 255 =>   sin_data_int <= to_unsigned(6246,N); cos_data_int <= to_unsigned(15146,N);
          when 256 =>   sin_data_int <= to_unsigned(6269,N); cos_data_int <= to_unsigned(15136,N);
          when 257 =>   sin_data_int <= to_unsigned(6293,N); cos_data_int <= to_unsigned(15127,N);
          when 258 =>   sin_data_int <= to_unsigned(6316,N); cos_data_int <= to_unsigned(15117,N);
          when 259 =>   sin_data_int <= to_unsigned(6339,N); cos_data_int <= to_unsigned(15107,N);
          when 260 =>   sin_data_int <= to_unsigned(6362,N); cos_data_int <= to_unsigned(15098,N);
          when 261 =>   sin_data_int <= to_unsigned(6385,N); cos_data_int <= to_unsigned(15088,N);
          when 262 =>   sin_data_int <= to_unsigned(6408,N); cos_data_int <= to_unsigned(15078,N);
          when 263 =>   sin_data_int <= to_unsigned(6432,N); cos_data_int <= to_unsigned(15068,N);
          when 264 =>   sin_data_int <= to_unsigned(6455,N); cos_data_int <= to_unsigned(15058,N);
          when 265 =>   sin_data_int <= to_unsigned(6478,N); cos_data_int <= to_unsigned(15048,N);
          when 266 =>   sin_data_int <= to_unsigned(6501,N); cos_data_int <= to_unsigned(15038,N);
          when 267 =>   sin_data_int <= to_unsigned(6524,N); cos_data_int <= to_unsigned(15028,N);
          when 268 =>   sin_data_int <= to_unsigned(6547,N); cos_data_int <= to_unsigned(15018,N);
          when 269 =>   sin_data_int <= to_unsigned(6570,N); cos_data_int <= to_unsigned(15008,N);
          when 270 =>   sin_data_int <= to_unsigned(6593,N); cos_data_int <= to_unsigned(14998,N);
          when 271 =>   sin_data_int <= to_unsigned(6616,N); cos_data_int <= to_unsigned(14988,N);
          when 272 =>   sin_data_int <= to_unsigned(6639,N); cos_data_int <= to_unsigned(14978,N);
          when 273 =>   sin_data_int <= to_unsigned(6662,N); cos_data_int <= to_unsigned(14968,N);
          when 274 =>   sin_data_int <= to_unsigned(6685,N); cos_data_int <= to_unsigned(14957,N);
          when 275 =>   sin_data_int <= to_unsigned(6708,N); cos_data_int <= to_unsigned(14947,N);
          when 276 =>   sin_data_int <= to_unsigned(6731,N); cos_data_int <= to_unsigned(14937,N);
          when 277 =>   sin_data_int <= to_unsigned(6754,N); cos_data_int <= to_unsigned(14927,N);
          when 278 =>   sin_data_int <= to_unsigned(6777,N); cos_data_int <= to_unsigned(14916,N);
          when 279 =>   sin_data_int <= to_unsigned(6799,N); cos_data_int <= to_unsigned(14906,N);
          when 280 =>   sin_data_int <= to_unsigned(6822,N); cos_data_int <= to_unsigned(14895,N);
          when 281 =>   sin_data_int <= to_unsigned(6845,N); cos_data_int <= to_unsigned(14885,N);
          when 282 =>   sin_data_int <= to_unsigned(6868,N); cos_data_int <= to_unsigned(14874,N);
          when 283 =>   sin_data_int <= to_unsigned(6891,N); cos_data_int <= to_unsigned(14864,N);
          when 284 =>   sin_data_int <= to_unsigned(6914,N); cos_data_int <= to_unsigned(14853,N);
          when 285 =>   sin_data_int <= to_unsigned(6936,N); cos_data_int <= to_unsigned(14843,N);
          when 286 =>   sin_data_int <= to_unsigned(6959,N); cos_data_int <= to_unsigned(14832,N);
          when 287 =>   sin_data_int <= to_unsigned(6982,N); cos_data_int <= to_unsigned(14821,N);
          when 288 =>   sin_data_int <= to_unsigned(7005,N); cos_data_int <= to_unsigned(14810,N);
          when 289 =>   sin_data_int <= to_unsigned(7027,N); cos_data_int <= to_unsigned(14800,N);
          when 290 =>   sin_data_int <= to_unsigned(7050,N); cos_data_int <= to_unsigned(14789,N);
          when 291 =>   sin_data_int <= to_unsigned(7073,N); cos_data_int <= to_unsigned(14778,N);
          when 292 =>   sin_data_int <= to_unsigned(7095,N); cos_data_int <= to_unsigned(14767,N);
          when 293 =>   sin_data_int <= to_unsigned(7118,N); cos_data_int <= to_unsigned(14756,N);
          when 294 =>   sin_data_int <= to_unsigned(7141,N); cos_data_int <= to_unsigned(14745,N);
          when 295 =>   sin_data_int <= to_unsigned(7163,N); cos_data_int <= to_unsigned(14734,N);
          when 296 =>   sin_data_int <= to_unsigned(7186,N); cos_data_int <= to_unsigned(14723,N);
          when 297 =>   sin_data_int <= to_unsigned(7208,N); cos_data_int <= to_unsigned(14712,N);
          when 298 =>   sin_data_int <= to_unsigned(7231,N); cos_data_int <= to_unsigned(14701,N);
          when 299 =>   sin_data_int <= to_unsigned(7253,N); cos_data_int <= to_unsigned(14690,N);
          when 300 =>   sin_data_int <= to_unsigned(7276,N); cos_data_int <= to_unsigned(14679,N);
          when 301 =>   sin_data_int <= to_unsigned(7299,N); cos_data_int <= to_unsigned(14668,N);
          when 302 =>   sin_data_int <= to_unsigned(7321,N); cos_data_int <= to_unsigned(14657,N);
          when 303 =>   sin_data_int <= to_unsigned(7343,N); cos_data_int <= to_unsigned(14645,N);
          when 304 =>   sin_data_int <= to_unsigned(7366,N); cos_data_int <= to_unsigned(14634,N);
          when 305 =>   sin_data_int <= to_unsigned(7388,N); cos_data_int <= to_unsigned(14623,N);
          when 306 =>   sin_data_int <= to_unsigned(7411,N); cos_data_int <= to_unsigned(14611,N);
          when 307 =>   sin_data_int <= to_unsigned(7433,N); cos_data_int <= to_unsigned(14600,N);
          when 308 =>   sin_data_int <= to_unsigned(7456,N); cos_data_int <= to_unsigned(14589,N);
          when 309 =>   sin_data_int <= to_unsigned(7478,N); cos_data_int <= to_unsigned(14577,N);
          when 310 =>   sin_data_int <= to_unsigned(7500,N); cos_data_int <= to_unsigned(14566,N);
          when 311 =>   sin_data_int <= to_unsigned(7523,N); cos_data_int <= to_unsigned(14554,N);
          when 312 =>   sin_data_int <= to_unsigned(7545,N); cos_data_int <= to_unsigned(14543,N);
          when 313 =>   sin_data_int <= to_unsigned(7567,N); cos_data_int <= to_unsigned(14531,N);
          when 314 =>   sin_data_int <= to_unsigned(7590,N); cos_data_int <= to_unsigned(14519,N);
          when 315 =>   sin_data_int <= to_unsigned(7612,N); cos_data_int <= to_unsigned(14508,N);
          when 316 =>   sin_data_int <= to_unsigned(7634,N); cos_data_int <= to_unsigned(14496,N);
          when 317 =>   sin_data_int <= to_unsigned(7656,N); cos_data_int <= to_unsigned(14484,N);
          when 318 =>   sin_data_int <= to_unsigned(7678,N); cos_data_int <= to_unsigned(14473,N);
          when 319 =>   sin_data_int <= to_unsigned(7701,N); cos_data_int <= to_unsigned(14461,N);
          when 320 =>   sin_data_int <= to_unsigned(7723,N); cos_data_int <= to_unsigned(14449,N);
          when 321 =>   sin_data_int <= to_unsigned(7745,N); cos_data_int <= to_unsigned(14437,N);
          when 322 =>   sin_data_int <= to_unsigned(7767,N); cos_data_int <= to_unsigned(14425,N);
          when 323 =>   sin_data_int <= to_unsigned(7789,N); cos_data_int <= to_unsigned(14413,N);
          when 324 =>   sin_data_int <= to_unsigned(7811,N); cos_data_int <= to_unsigned(14401,N);
          when 325 =>   sin_data_int <= to_unsigned(7833,N); cos_data_int <= to_unsigned(14389,N);
          when 326 =>   sin_data_int <= to_unsigned(7856,N); cos_data_int <= to_unsigned(14377,N);
          when 327 =>   sin_data_int <= to_unsigned(7878,N); cos_data_int <= to_unsigned(14365,N);
          when 328 =>   sin_data_int <= to_unsigned(7900,N); cos_data_int <= to_unsigned(14353,N);
          when 329 =>   sin_data_int <= to_unsigned(7922,N); cos_data_int <= to_unsigned(14341,N);
          when 330 =>   sin_data_int <= to_unsigned(7944,N); cos_data_int <= to_unsigned(14329,N);
          when 331 =>   sin_data_int <= to_unsigned(7966,N); cos_data_int <= to_unsigned(14317,N);
          when 332 =>   sin_data_int <= to_unsigned(7988,N); cos_data_int <= to_unsigned(14304,N);
          when 333 =>   sin_data_int <= to_unsigned(8009,N); cos_data_int <= to_unsigned(14292,N);
          when 334 =>   sin_data_int <= to_unsigned(8031,N); cos_data_int <= to_unsigned(14280,N);
          when 335 =>   sin_data_int <= to_unsigned(8053,N); cos_data_int <= to_unsigned(14267,N);
          when 336 =>   sin_data_int <= to_unsigned(8075,N); cos_data_int <= to_unsigned(14255,N);
          when 337 =>   sin_data_int <= to_unsigned(8097,N); cos_data_int <= to_unsigned(14243,N);
          when 338 =>   sin_data_int <= to_unsigned(8119,N); cos_data_int <= to_unsigned(14230,N);
          when 339 =>   sin_data_int <= to_unsigned(8141,N); cos_data_int <= to_unsigned(14218,N);
          when 340 =>   sin_data_int <= to_unsigned(8162,N); cos_data_int <= to_unsigned(14205,N);
          when 341 =>   sin_data_int <= to_unsigned(8184,N); cos_data_int <= to_unsigned(14193,N);
          when 342 =>   sin_data_int <= to_unsigned(8206,N); cos_data_int <= to_unsigned(14180,N);
          when 343 =>   sin_data_int <= to_unsigned(8228,N); cos_data_int <= to_unsigned(14167,N);
          when 344 =>   sin_data_int <= to_unsigned(8249,N); cos_data_int <= to_unsigned(14155,N);
          when 345 =>   sin_data_int <= to_unsigned(8271,N); cos_data_int <= to_unsigned(14142,N);
          when 346 =>   sin_data_int <= to_unsigned(8293,N); cos_data_int <= to_unsigned(14129,N);
          when 347 =>   sin_data_int <= to_unsigned(8315,N); cos_data_int <= to_unsigned(14117,N);
          when 348 =>   sin_data_int <= to_unsigned(8336,N); cos_data_int <= to_unsigned(14104,N);
          when 349 =>   sin_data_int <= to_unsigned(8358,N); cos_data_int <= to_unsigned(14091,N);
          when 350 =>   sin_data_int <= to_unsigned(8379,N); cos_data_int <= to_unsigned(14078,N);
          when 351 =>   sin_data_int <= to_unsigned(8401,N); cos_data_int <= to_unsigned(14065,N);
          when 352 =>   sin_data_int <= to_unsigned(8423,N); cos_data_int <= to_unsigned(14053,N);
          when 353 =>   sin_data_int <= to_unsigned(8444,N); cos_data_int <= to_unsigned(14040,N);
          when 354 =>   sin_data_int <= to_unsigned(8466,N); cos_data_int <= to_unsigned(14027,N);
          when 355 =>   sin_data_int <= to_unsigned(8487,N); cos_data_int <= to_unsigned(14014,N);
          when 356 =>   sin_data_int <= to_unsigned(8509,N); cos_data_int <= to_unsigned(14001,N);
          when 357 =>   sin_data_int <= to_unsigned(8530,N); cos_data_int <= to_unsigned(13988,N);
          when 358 =>   sin_data_int <= to_unsigned(8552,N); cos_data_int <= to_unsigned(13974,N);
          when 359 =>   sin_data_int <= to_unsigned(8573,N); cos_data_int <= to_unsigned(13961,N);
          when 360 =>   sin_data_int <= to_unsigned(8594,N); cos_data_int <= to_unsigned(13948,N);
          when 361 =>   sin_data_int <= to_unsigned(8616,N); cos_data_int <= to_unsigned(13935,N);
          when 362 =>   sin_data_int <= to_unsigned(8637,N); cos_data_int <= to_unsigned(13922,N);
          when 363 =>   sin_data_int <= to_unsigned(8658,N); cos_data_int <= to_unsigned(13908,N);
          when 364 =>   sin_data_int <= to_unsigned(8680,N); cos_data_int <= to_unsigned(13895,N);
          when 365 =>   sin_data_int <= to_unsigned(8701,N); cos_data_int <= to_unsigned(13882,N);
          when 366 =>   sin_data_int <= to_unsigned(8722,N); cos_data_int <= to_unsigned(13868,N);
          when 367 =>   sin_data_int <= to_unsigned(8744,N); cos_data_int <= to_unsigned(13855,N);
          when 368 =>   sin_data_int <= to_unsigned(8765,N); cos_data_int <= to_unsigned(13842,N);
          when 369 =>   sin_data_int <= to_unsigned(8786,N); cos_data_int <= to_unsigned(13828,N);
          when 370 =>   sin_data_int <= to_unsigned(8807,N); cos_data_int <= to_unsigned(13815,N);
          when 371 =>   sin_data_int <= to_unsigned(8829,N); cos_data_int <= to_unsigned(13801,N);
          when 372 =>   sin_data_int <= to_unsigned(8850,N); cos_data_int <= to_unsigned(13788,N);
          when 373 =>   sin_data_int <= to_unsigned(8871,N); cos_data_int <= to_unsigned(13774,N);
          when 374 =>   sin_data_int <= to_unsigned(8892,N); cos_data_int <= to_unsigned(13760,N);
          when 375 =>   sin_data_int <= to_unsigned(8913,N); cos_data_int <= to_unsigned(13747,N);
          when 376 =>   sin_data_int <= to_unsigned(8934,N); cos_data_int <= to_unsigned(13733,N);
          when 377 =>   sin_data_int <= to_unsigned(8955,N); cos_data_int <= to_unsigned(13719,N);
          when 378 =>   sin_data_int <= to_unsigned(8976,N); cos_data_int <= to_unsigned(13705,N);
          when 379 =>   sin_data_int <= to_unsigned(8997,N); cos_data_int <= to_unsigned(13692,N);
          when 380 =>   sin_data_int <= to_unsigned(9018,N); cos_data_int <= to_unsigned(13678,N);
          when 381 =>   sin_data_int <= to_unsigned(9039,N); cos_data_int <= to_unsigned(13664,N);
          when 382 =>   sin_data_int <= to_unsigned(9060,N); cos_data_int <= to_unsigned(13650,N);
          when 383 =>   sin_data_int <= to_unsigned(9081,N); cos_data_int <= to_unsigned(13636,N);
          when 384 =>   sin_data_int <= to_unsigned(9102,N); cos_data_int <= to_unsigned(13622,N);
          when 385 =>   sin_data_int <= to_unsigned(9123,N); cos_data_int <= to_unsigned(13608,N);
          when 386 =>   sin_data_int <= to_unsigned(9144,N); cos_data_int <= to_unsigned(13594,N);
          when 387 =>   sin_data_int <= to_unsigned(9165,N); cos_data_int <= to_unsigned(13580,N);
          when 388 =>   sin_data_int <= to_unsigned(9185,N); cos_data_int <= to_unsigned(13566,N);
          when 389 =>   sin_data_int <= to_unsigned(9206,N); cos_data_int <= to_unsigned(13552,N);
          when 390 =>   sin_data_int <= to_unsigned(9227,N); cos_data_int <= to_unsigned(13538,N);
          when 391 =>   sin_data_int <= to_unsigned(9248,N); cos_data_int <= to_unsigned(13524,N);
          when 392 =>   sin_data_int <= to_unsigned(9268,N); cos_data_int <= to_unsigned(13510,N);
          when 393 =>   sin_data_int <= to_unsigned(9289,N); cos_data_int <= to_unsigned(13495,N);
          when 394 =>   sin_data_int <= to_unsigned(9310,N); cos_data_int <= to_unsigned(13481,N);
          when 395 =>   sin_data_int <= to_unsigned(9331,N); cos_data_int <= to_unsigned(13467,N);
          when 396 =>   sin_data_int <= to_unsigned(9351,N); cos_data_int <= to_unsigned(13452,N);
          when 397 =>   sin_data_int <= to_unsigned(9372,N); cos_data_int <= to_unsigned(13438,N);
          when 398 =>   sin_data_int <= to_unsigned(9392,N); cos_data_int <= to_unsigned(13424,N);
          when 399 =>   sin_data_int <= to_unsigned(9413,N); cos_data_int <= to_unsigned(13409,N);
          when 400 =>   sin_data_int <= to_unsigned(9434,N); cos_data_int <= to_unsigned(13395,N);
          when 401 =>   sin_data_int <= to_unsigned(9454,N); cos_data_int <= to_unsigned(13380,N);
          when 402 =>   sin_data_int <= to_unsigned(9475,N); cos_data_int <= to_unsigned(13366,N);
          when 403 =>   sin_data_int <= to_unsigned(9495,N); cos_data_int <= to_unsigned(13351,N);
          when 404 =>   sin_data_int <= to_unsigned(9516,N); cos_data_int <= to_unsigned(13337,N);
          when 405 =>   sin_data_int <= to_unsigned(9536,N); cos_data_int <= to_unsigned(13322,N);
          when 406 =>   sin_data_int <= to_unsigned(9556,N); cos_data_int <= to_unsigned(13307,N);
          when 407 =>   sin_data_int <= to_unsigned(9577,N); cos_data_int <= to_unsigned(13293,N);
          when 408 =>   sin_data_int <= to_unsigned(9597,N); cos_data_int <= to_unsigned(13278,N);
          when 409 =>   sin_data_int <= to_unsigned(9618,N); cos_data_int <= to_unsigned(13263,N);
          when 410 =>   sin_data_int <= to_unsigned(9638,N); cos_data_int <= to_unsigned(13249,N);
          when 411 =>   sin_data_int <= to_unsigned(9658,N); cos_data_int <= to_unsigned(13234,N);
          when 412 =>   sin_data_int <= to_unsigned(9679,N); cos_data_int <= to_unsigned(13219,N);
          when 413 =>   sin_data_int <= to_unsigned(9699,N); cos_data_int <= to_unsigned(13204,N);
          when 414 =>   sin_data_int <= to_unsigned(9719,N); cos_data_int <= to_unsigned(13189,N);
          when 415 =>   sin_data_int <= to_unsigned(9739,N); cos_data_int <= to_unsigned(13174,N);
          when 416 =>   sin_data_int <= to_unsigned(9759,N); cos_data_int <= to_unsigned(13159,N);
          when 417 =>   sin_data_int <= to_unsigned(9780,N); cos_data_int <= to_unsigned(13144,N);
          when 418 =>   sin_data_int <= to_unsigned(9800,N); cos_data_int <= to_unsigned(13129,N);
          when 419 =>   sin_data_int <= to_unsigned(9820,N); cos_data_int <= to_unsigned(13114,N);
          when 420 =>   sin_data_int <= to_unsigned(9840,N); cos_data_int <= to_unsigned(13099,N);
          when 421 =>   sin_data_int <= to_unsigned(9860,N); cos_data_int <= to_unsigned(13084,N);
          when 422 =>   sin_data_int <= to_unsigned(9880,N); cos_data_int <= to_unsigned(13069,N);
          when 423 =>   sin_data_int <= to_unsigned(9900,N); cos_data_int <= to_unsigned(13054,N);
          when 424 =>   sin_data_int <= to_unsigned(9920,N); cos_data_int <= to_unsigned(13038,N);
          when 425 =>   sin_data_int <= to_unsigned(9940,N); cos_data_int <= to_unsigned(13023,N);
          when 426 =>   sin_data_int <= to_unsigned(9960,N); cos_data_int <= to_unsigned(13008,N);
          when 427 =>   sin_data_int <= to_unsigned(9980,N); cos_data_int <= to_unsigned(12993,N);
          when 428 =>   sin_data_int <= to_unsigned(10000,N); cos_data_int <= to_unsigned(12977,N);
          when 429 =>   sin_data_int <= to_unsigned(10020,N); cos_data_int <= to_unsigned(12962,N);
          when 430 =>   sin_data_int <= to_unsigned(10040,N); cos_data_int <= to_unsigned(12947,N);
          when 431 =>   sin_data_int <= to_unsigned(10060,N); cos_data_int <= to_unsigned(12931,N);
          when 432 =>   sin_data_int <= to_unsigned(10079,N); cos_data_int <= to_unsigned(12916,N);
          when 433 =>   sin_data_int <= to_unsigned(10099,N); cos_data_int <= to_unsigned(12900,N);
          when 434 =>   sin_data_int <= to_unsigned(10119,N); cos_data_int <= to_unsigned(12885,N);
          when 435 =>   sin_data_int <= to_unsigned(10139,N); cos_data_int <= to_unsigned(12869,N);
          when 436 =>   sin_data_int <= to_unsigned(10159,N); cos_data_int <= to_unsigned(12854,N);
          when 437 =>   sin_data_int <= to_unsigned(10178,N); cos_data_int <= to_unsigned(12838,N);
          when 438 =>   sin_data_int <= to_unsigned(10198,N); cos_data_int <= to_unsigned(12822,N);
          when 439 =>   sin_data_int <= to_unsigned(10218,N); cos_data_int <= to_unsigned(12807,N);
          when 440 =>   sin_data_int <= to_unsigned(10237,N); cos_data_int <= to_unsigned(12791,N);
          when 441 =>   sin_data_int <= to_unsigned(10257,N); cos_data_int <= to_unsigned(12775,N);
          when 442 =>   sin_data_int <= to_unsigned(10276,N); cos_data_int <= to_unsigned(12760,N);
          when 443 =>   sin_data_int <= to_unsigned(10296,N); cos_data_int <= to_unsigned(12744,N);
          when 444 =>   sin_data_int <= to_unsigned(10315,N); cos_data_int <= to_unsigned(12728,N);
          when 445 =>   sin_data_int <= to_unsigned(10335,N); cos_data_int <= to_unsigned(12712,N);
          when 446 =>   sin_data_int <= to_unsigned(10354,N); cos_data_int <= to_unsigned(12696,N);
          when 447 =>   sin_data_int <= to_unsigned(10374,N); cos_data_int <= to_unsigned(12680,N);
          when 448 =>   sin_data_int <= to_unsigned(10393,N); cos_data_int <= to_unsigned(12665,N);
          when 449 =>   sin_data_int <= to_unsigned(10413,N); cos_data_int <= to_unsigned(12649,N);
          when 450 =>   sin_data_int <= to_unsigned(10432,N); cos_data_int <= to_unsigned(12633,N);
          when 451 =>   sin_data_int <= to_unsigned(10452,N); cos_data_int <= to_unsigned(12617,N);
          when 452 =>   sin_data_int <= to_unsigned(10471,N); cos_data_int <= to_unsigned(12600,N);
          when 453 =>   sin_data_int <= to_unsigned(10490,N); cos_data_int <= to_unsigned(12584,N);
          when 454 =>   sin_data_int <= to_unsigned(10510,N); cos_data_int <= to_unsigned(12568,N);
          when 455 =>   sin_data_int <= to_unsigned(10529,N); cos_data_int <= to_unsigned(12552,N);
          when 456 =>   sin_data_int <= to_unsigned(10548,N); cos_data_int <= to_unsigned(12536,N);
          when 457 =>   sin_data_int <= to_unsigned(10567,N); cos_data_int <= to_unsigned(12520,N);
          when 458 =>   sin_data_int <= to_unsigned(10586,N); cos_data_int <= to_unsigned(12504,N);
          when 459 =>   sin_data_int <= to_unsigned(10606,N); cos_data_int <= to_unsigned(12487,N);
          when 460 =>   sin_data_int <= to_unsigned(10625,N); cos_data_int <= to_unsigned(12471,N);
          when 461 =>   sin_data_int <= to_unsigned(10644,N); cos_data_int <= to_unsigned(12455,N);
          when 462 =>   sin_data_int <= to_unsigned(10663,N); cos_data_int <= to_unsigned(12438,N);
          when 463 =>   sin_data_int <= to_unsigned(10682,N); cos_data_int <= to_unsigned(12422,N);
          when 464 =>   sin_data_int <= to_unsigned(10701,N); cos_data_int <= to_unsigned(12406,N);
          when 465 =>   sin_data_int <= to_unsigned(10720,N); cos_data_int <= to_unsigned(12389,N);
          when 466 =>   sin_data_int <= to_unsigned(10739,N); cos_data_int <= to_unsigned(12373,N);
          when 467 =>   sin_data_int <= to_unsigned(10758,N); cos_data_int <= to_unsigned(12356,N);
          when 468 =>   sin_data_int <= to_unsigned(10777,N); cos_data_int <= to_unsigned(12340,N);
          when 469 =>   sin_data_int <= to_unsigned(10796,N); cos_data_int <= to_unsigned(12323,N);
          when 470 =>   sin_data_int <= to_unsigned(10815,N); cos_data_int <= to_unsigned(12307,N);
          when 471 =>   sin_data_int <= to_unsigned(10834,N); cos_data_int <= to_unsigned(12290,N);
          when 472 =>   sin_data_int <= to_unsigned(10853,N); cos_data_int <= to_unsigned(12273,N);
          when 473 =>   sin_data_int <= to_unsigned(10871,N); cos_data_int <= to_unsigned(12257,N);
          when 474 =>   sin_data_int <= to_unsigned(10890,N); cos_data_int <= to_unsigned(12240,N);
          when 475 =>   sin_data_int <= to_unsigned(10909,N); cos_data_int <= to_unsigned(12223,N);
          when 476 =>   sin_data_int <= to_unsigned(10928,N); cos_data_int <= to_unsigned(12207,N);
          when 477 =>   sin_data_int <= to_unsigned(10946,N); cos_data_int <= to_unsigned(12190,N);
          when 478 =>   sin_data_int <= to_unsigned(10965,N); cos_data_int <= to_unsigned(12173,N);
          when 479 =>   sin_data_int <= to_unsigned(10984,N); cos_data_int <= to_unsigned(12156,N);
          when 480 =>   sin_data_int <= to_unsigned(11002,N); cos_data_int <= to_unsigned(12139,N);
          when 481 =>   sin_data_int <= to_unsigned(11021,N); cos_data_int <= to_unsigned(12122,N);
          when 482 =>   sin_data_int <= to_unsigned(11040,N); cos_data_int <= to_unsigned(12105,N);
          when 483 =>   sin_data_int <= to_unsigned(11058,N); cos_data_int <= to_unsigned(12088,N);
          when 484 =>   sin_data_int <= to_unsigned(11077,N); cos_data_int <= to_unsigned(12072,N);
          when 485 =>   sin_data_int <= to_unsigned(11095,N); cos_data_int <= to_unsigned(12054,N);
          when 486 =>   sin_data_int <= to_unsigned(11114,N); cos_data_int <= to_unsigned(12037,N);
          when 487 =>   sin_data_int <= to_unsigned(11132,N); cos_data_int <= to_unsigned(12020,N);
          when 488 =>   sin_data_int <= to_unsigned(11150,N); cos_data_int <= to_unsigned(12003,N);
          when 489 =>   sin_data_int <= to_unsigned(11169,N); cos_data_int <= to_unsigned(11986,N);
          when 490 =>   sin_data_int <= to_unsigned(11187,N); cos_data_int <= to_unsigned(11969,N);
          when 491 =>   sin_data_int <= to_unsigned(11206,N); cos_data_int <= to_unsigned(11952,N);
          when 492 =>   sin_data_int <= to_unsigned(11224,N); cos_data_int <= to_unsigned(11935,N);
          when 493 =>   sin_data_int <= to_unsigned(11242,N); cos_data_int <= to_unsigned(11917,N);
          when 494 =>   sin_data_int <= to_unsigned(11260,N); cos_data_int <= to_unsigned(11900,N);
          when 495 =>   sin_data_int <= to_unsigned(11279,N); cos_data_int <= to_unsigned(11883,N);
          when 496 =>   sin_data_int <= to_unsigned(11297,N); cos_data_int <= to_unsigned(11866,N);
          when 497 =>   sin_data_int <= to_unsigned(11315,N); cos_data_int <= to_unsigned(11848,N);
          when 498 =>   sin_data_int <= to_unsigned(11333,N); cos_data_int <= to_unsigned(11831,N);
          when 499 =>   sin_data_int <= to_unsigned(11351,N); cos_data_int <= to_unsigned(11813,N);
          when 500 =>   sin_data_int <= to_unsigned(11370,N); cos_data_int <= to_unsigned(11796,N);
          when 501 =>   sin_data_int <= to_unsigned(11388,N); cos_data_int <= to_unsigned(11779,N);
          when 502 =>   sin_data_int <= to_unsigned(11406,N); cos_data_int <= to_unsigned(11761,N);
          when 503 =>   sin_data_int <= to_unsigned(11424,N); cos_data_int <= to_unsigned(11744,N);
          when 504 =>   sin_data_int <= to_unsigned(11442,N); cos_data_int <= to_unsigned(11726,N);
          when 505 =>   sin_data_int <= to_unsigned(11460,N); cos_data_int <= to_unsigned(11708,N);
          when 506 =>   sin_data_int <= to_unsigned(11478,N); cos_data_int <= to_unsigned(11691,N);
          when 507 =>   sin_data_int <= to_unsigned(11496,N); cos_data_int <= to_unsigned(11673,N);
          when 508 =>   sin_data_int <= to_unsigned(11513,N); cos_data_int <= to_unsigned(11656,N);
          when 509 =>   sin_data_int <= to_unsigned(11531,N); cos_data_int <= to_unsigned(11638,N);
          when 510 =>   sin_data_int <= to_unsigned(11549,N); cos_data_int <= to_unsigned(11620,N);
          when 511 =>   sin_data_int <= to_unsigned(11567,N); cos_data_int <= to_unsigned(11602,N);
          when 512 =>   sin_data_int <= to_unsigned(11585,N); cos_data_int <= to_unsigned(11585,N);
          when 513 =>   sin_data_int <= to_unsigned(11602,N); cos_data_int <= to_unsigned(11567,N);
          when 514 =>   sin_data_int <= to_unsigned(11620,N); cos_data_int <= to_unsigned(11549,N);
          when 515 =>   sin_data_int <= to_unsigned(11638,N); cos_data_int <= to_unsigned(11531,N);
          when 516 =>   sin_data_int <= to_unsigned(11656,N); cos_data_int <= to_unsigned(11513,N);
          when 517 =>   sin_data_int <= to_unsigned(11673,N); cos_data_int <= to_unsigned(11496,N);
          when 518 =>   sin_data_int <= to_unsigned(11691,N); cos_data_int <= to_unsigned(11478,N);
          when 519 =>   sin_data_int <= to_unsigned(11708,N); cos_data_int <= to_unsigned(11460,N);
          when 520 =>   sin_data_int <= to_unsigned(11726,N); cos_data_int <= to_unsigned(11442,N);
          when 521 =>   sin_data_int <= to_unsigned(11744,N); cos_data_int <= to_unsigned(11424,N);
          when 522 =>   sin_data_int <= to_unsigned(11761,N); cos_data_int <= to_unsigned(11406,N);
          when 523 =>   sin_data_int <= to_unsigned(11779,N); cos_data_int <= to_unsigned(11388,N);
          when 524 =>   sin_data_int <= to_unsigned(11796,N); cos_data_int <= to_unsigned(11370,N);
          when 525 =>   sin_data_int <= to_unsigned(11813,N); cos_data_int <= to_unsigned(11351,N);
          when 526 =>   sin_data_int <= to_unsigned(11831,N); cos_data_int <= to_unsigned(11333,N);
          when 527 =>   sin_data_int <= to_unsigned(11848,N); cos_data_int <= to_unsigned(11315,N);
          when 528 =>   sin_data_int <= to_unsigned(11866,N); cos_data_int <= to_unsigned(11297,N);
          when 529 =>   sin_data_int <= to_unsigned(11883,N); cos_data_int <= to_unsigned(11279,N);
          when 530 =>   sin_data_int <= to_unsigned(11900,N); cos_data_int <= to_unsigned(11260,N);
          when 531 =>   sin_data_int <= to_unsigned(11917,N); cos_data_int <= to_unsigned(11242,N);
          when 532 =>   sin_data_int <= to_unsigned(11935,N); cos_data_int <= to_unsigned(11224,N);
          when 533 =>   sin_data_int <= to_unsigned(11952,N); cos_data_int <= to_unsigned(11206,N);
          when 534 =>   sin_data_int <= to_unsigned(11969,N); cos_data_int <= to_unsigned(11187,N);
          when 535 =>   sin_data_int <= to_unsigned(11986,N); cos_data_int <= to_unsigned(11169,N);
          when 536 =>   sin_data_int <= to_unsigned(12003,N); cos_data_int <= to_unsigned(11150,N);
          when 537 =>   sin_data_int <= to_unsigned(12020,N); cos_data_int <= to_unsigned(11132,N);
          when 538 =>   sin_data_int <= to_unsigned(12037,N); cos_data_int <= to_unsigned(11114,N);
          when 539 =>   sin_data_int <= to_unsigned(12054,N); cos_data_int <= to_unsigned(11095,N);
          when 540 =>   sin_data_int <= to_unsigned(12072,N); cos_data_int <= to_unsigned(11077,N);
          when 541 =>   sin_data_int <= to_unsigned(12088,N); cos_data_int <= to_unsigned(11058,N);
          when 542 =>   sin_data_int <= to_unsigned(12105,N); cos_data_int <= to_unsigned(11040,N);
          when 543 =>   sin_data_int <= to_unsigned(12122,N); cos_data_int <= to_unsigned(11021,N);
          when 544 =>   sin_data_int <= to_unsigned(12139,N); cos_data_int <= to_unsigned(11002,N);
          when 545 =>   sin_data_int <= to_unsigned(12156,N); cos_data_int <= to_unsigned(10984,N);
          when 546 =>   sin_data_int <= to_unsigned(12173,N); cos_data_int <= to_unsigned(10965,N);
          when 547 =>   sin_data_int <= to_unsigned(12190,N); cos_data_int <= to_unsigned(10946,N);
          when 548 =>   sin_data_int <= to_unsigned(12207,N); cos_data_int <= to_unsigned(10928,N);
          when 549 =>   sin_data_int <= to_unsigned(12223,N); cos_data_int <= to_unsigned(10909,N);
          when 550 =>   sin_data_int <= to_unsigned(12240,N); cos_data_int <= to_unsigned(10890,N);
          when 551 =>   sin_data_int <= to_unsigned(12257,N); cos_data_int <= to_unsigned(10871,N);
          when 552 =>   sin_data_int <= to_unsigned(12273,N); cos_data_int <= to_unsigned(10853,N);
          when 553 =>   sin_data_int <= to_unsigned(12290,N); cos_data_int <= to_unsigned(10834,N);
          when 554 =>   sin_data_int <= to_unsigned(12307,N); cos_data_int <= to_unsigned(10815,N);
          when 555 =>   sin_data_int <= to_unsigned(12323,N); cos_data_int <= to_unsigned(10796,N);
          when 556 =>   sin_data_int <= to_unsigned(12340,N); cos_data_int <= to_unsigned(10777,N);
          when 557 =>   sin_data_int <= to_unsigned(12356,N); cos_data_int <= to_unsigned(10758,N);
          when 558 =>   sin_data_int <= to_unsigned(12373,N); cos_data_int <= to_unsigned(10739,N);
          when 559 =>   sin_data_int <= to_unsigned(12389,N); cos_data_int <= to_unsigned(10720,N);
          when 560 =>   sin_data_int <= to_unsigned(12406,N); cos_data_int <= to_unsigned(10701,N);
          when 561 =>   sin_data_int <= to_unsigned(12422,N); cos_data_int <= to_unsigned(10682,N);
          when 562 =>   sin_data_int <= to_unsigned(12438,N); cos_data_int <= to_unsigned(10663,N);
          when 563 =>   sin_data_int <= to_unsigned(12455,N); cos_data_int <= to_unsigned(10644,N);
          when 564 =>   sin_data_int <= to_unsigned(12471,N); cos_data_int <= to_unsigned(10625,N);
          when 565 =>   sin_data_int <= to_unsigned(12487,N); cos_data_int <= to_unsigned(10606,N);
          when 566 =>   sin_data_int <= to_unsigned(12504,N); cos_data_int <= to_unsigned(10586,N);
          when 567 =>   sin_data_int <= to_unsigned(12520,N); cos_data_int <= to_unsigned(10567,N);
          when 568 =>   sin_data_int <= to_unsigned(12536,N); cos_data_int <= to_unsigned(10548,N);
          when 569 =>   sin_data_int <= to_unsigned(12552,N); cos_data_int <= to_unsigned(10529,N);
          when 570 =>   sin_data_int <= to_unsigned(12568,N); cos_data_int <= to_unsigned(10510,N);
          when 571 =>   sin_data_int <= to_unsigned(12584,N); cos_data_int <= to_unsigned(10490,N);
          when 572 =>   sin_data_int <= to_unsigned(12600,N); cos_data_int <= to_unsigned(10471,N);
          when 573 =>   sin_data_int <= to_unsigned(12617,N); cos_data_int <= to_unsigned(10452,N);
          when 574 =>   sin_data_int <= to_unsigned(12633,N); cos_data_int <= to_unsigned(10432,N);
          when 575 =>   sin_data_int <= to_unsigned(12649,N); cos_data_int <= to_unsigned(10413,N);
          when 576 =>   sin_data_int <= to_unsigned(12665,N); cos_data_int <= to_unsigned(10393,N);
          when 577 =>   sin_data_int <= to_unsigned(12680,N); cos_data_int <= to_unsigned(10374,N);
          when 578 =>   sin_data_int <= to_unsigned(12696,N); cos_data_int <= to_unsigned(10354,N);
          when 579 =>   sin_data_int <= to_unsigned(12712,N); cos_data_int <= to_unsigned(10335,N);
          when 580 =>   sin_data_int <= to_unsigned(12728,N); cos_data_int <= to_unsigned(10315,N);
          when 581 =>   sin_data_int <= to_unsigned(12744,N); cos_data_int <= to_unsigned(10296,N);
          when 582 =>   sin_data_int <= to_unsigned(12760,N); cos_data_int <= to_unsigned(10276,N);
          when 583 =>   sin_data_int <= to_unsigned(12775,N); cos_data_int <= to_unsigned(10257,N);
          when 584 =>   sin_data_int <= to_unsigned(12791,N); cos_data_int <= to_unsigned(10237,N);
          when 585 =>   sin_data_int <= to_unsigned(12807,N); cos_data_int <= to_unsigned(10218,N);
          when 586 =>   sin_data_int <= to_unsigned(12822,N); cos_data_int <= to_unsigned(10198,N);
          when 587 =>   sin_data_int <= to_unsigned(12838,N); cos_data_int <= to_unsigned(10178,N);
          when 588 =>   sin_data_int <= to_unsigned(12854,N); cos_data_int <= to_unsigned(10159,N);
          when 589 =>   sin_data_int <= to_unsigned(12869,N); cos_data_int <= to_unsigned(10139,N);
          when 590 =>   sin_data_int <= to_unsigned(12885,N); cos_data_int <= to_unsigned(10119,N);
          when 591 =>   sin_data_int <= to_unsigned(12900,N); cos_data_int <= to_unsigned(10099,N);
          when 592 =>   sin_data_int <= to_unsigned(12916,N); cos_data_int <= to_unsigned(10079,N);
          when 593 =>   sin_data_int <= to_unsigned(12931,N); cos_data_int <= to_unsigned(10060,N);
          when 594 =>   sin_data_int <= to_unsigned(12947,N); cos_data_int <= to_unsigned(10040,N);
          when 595 =>   sin_data_int <= to_unsigned(12962,N); cos_data_int <= to_unsigned(10020,N);
          when 596 =>   sin_data_int <= to_unsigned(12977,N); cos_data_int <= to_unsigned(10000,N);
          when 597 =>   sin_data_int <= to_unsigned(12993,N); cos_data_int <= to_unsigned(9980,N);
          when 598 =>   sin_data_int <= to_unsigned(13008,N); cos_data_int <= to_unsigned(9960,N);
          when 599 =>   sin_data_int <= to_unsigned(13023,N); cos_data_int <= to_unsigned(9940,N);
          when 600 =>   sin_data_int <= to_unsigned(13038,N); cos_data_int <= to_unsigned(9920,N);
          when 601 =>   sin_data_int <= to_unsigned(13054,N); cos_data_int <= to_unsigned(9900,N);
          when 602 =>   sin_data_int <= to_unsigned(13069,N); cos_data_int <= to_unsigned(9880,N);
          when 603 =>   sin_data_int <= to_unsigned(13084,N); cos_data_int <= to_unsigned(9860,N);
          when 604 =>   sin_data_int <= to_unsigned(13099,N); cos_data_int <= to_unsigned(9840,N);
          when 605 =>   sin_data_int <= to_unsigned(13114,N); cos_data_int <= to_unsigned(9820,N);
          when 606 =>   sin_data_int <= to_unsigned(13129,N); cos_data_int <= to_unsigned(9800,N);
          when 607 =>   sin_data_int <= to_unsigned(13144,N); cos_data_int <= to_unsigned(9780,N);
          when 608 =>   sin_data_int <= to_unsigned(13159,N); cos_data_int <= to_unsigned(9759,N);
          when 609 =>   sin_data_int <= to_unsigned(13174,N); cos_data_int <= to_unsigned(9739,N);
          when 610 =>   sin_data_int <= to_unsigned(13189,N); cos_data_int <= to_unsigned(9719,N);
          when 611 =>   sin_data_int <= to_unsigned(13204,N); cos_data_int <= to_unsigned(9699,N);
          when 612 =>   sin_data_int <= to_unsigned(13219,N); cos_data_int <= to_unsigned(9679,N);
          when 613 =>   sin_data_int <= to_unsigned(13234,N); cos_data_int <= to_unsigned(9658,N);
          when 614 =>   sin_data_int <= to_unsigned(13249,N); cos_data_int <= to_unsigned(9638,N);
          when 615 =>   sin_data_int <= to_unsigned(13263,N); cos_data_int <= to_unsigned(9618,N);
          when 616 =>   sin_data_int <= to_unsigned(13278,N); cos_data_int <= to_unsigned(9597,N);
          when 617 =>   sin_data_int <= to_unsigned(13293,N); cos_data_int <= to_unsigned(9577,N);
          when 618 =>   sin_data_int <= to_unsigned(13307,N); cos_data_int <= to_unsigned(9556,N);
          when 619 =>   sin_data_int <= to_unsigned(13322,N); cos_data_int <= to_unsigned(9536,N);
          when 620 =>   sin_data_int <= to_unsigned(13337,N); cos_data_int <= to_unsigned(9516,N);
          when 621 =>   sin_data_int <= to_unsigned(13351,N); cos_data_int <= to_unsigned(9495,N);
          when 622 =>   sin_data_int <= to_unsigned(13366,N); cos_data_int <= to_unsigned(9475,N);
          when 623 =>   sin_data_int <= to_unsigned(13380,N); cos_data_int <= to_unsigned(9454,N);
          when 624 =>   sin_data_int <= to_unsigned(13395,N); cos_data_int <= to_unsigned(9434,N);
          when 625 =>   sin_data_int <= to_unsigned(13409,N); cos_data_int <= to_unsigned(9413,N);
          when 626 =>   sin_data_int <= to_unsigned(13424,N); cos_data_int <= to_unsigned(9392,N);
          when 627 =>   sin_data_int <= to_unsigned(13438,N); cos_data_int <= to_unsigned(9372,N);
          when 628 =>   sin_data_int <= to_unsigned(13452,N); cos_data_int <= to_unsigned(9351,N);
          when 629 =>   sin_data_int <= to_unsigned(13467,N); cos_data_int <= to_unsigned(9331,N);
          when 630 =>   sin_data_int <= to_unsigned(13481,N); cos_data_int <= to_unsigned(9310,N);
          when 631 =>   sin_data_int <= to_unsigned(13495,N); cos_data_int <= to_unsigned(9289,N);
          when 632 =>   sin_data_int <= to_unsigned(13510,N); cos_data_int <= to_unsigned(9268,N);
          when 633 =>   sin_data_int <= to_unsigned(13524,N); cos_data_int <= to_unsigned(9248,N);
          when 634 =>   sin_data_int <= to_unsigned(13538,N); cos_data_int <= to_unsigned(9227,N);
          when 635 =>   sin_data_int <= to_unsigned(13552,N); cos_data_int <= to_unsigned(9206,N);
          when 636 =>   sin_data_int <= to_unsigned(13566,N); cos_data_int <= to_unsigned(9185,N);
          when 637 =>   sin_data_int <= to_unsigned(13580,N); cos_data_int <= to_unsigned(9165,N);
          when 638 =>   sin_data_int <= to_unsigned(13594,N); cos_data_int <= to_unsigned(9144,N);
          when 639 =>   sin_data_int <= to_unsigned(13608,N); cos_data_int <= to_unsigned(9123,N);
          when 640 =>   sin_data_int <= to_unsigned(13622,N); cos_data_int <= to_unsigned(9102,N);
          when 641 =>   sin_data_int <= to_unsigned(13636,N); cos_data_int <= to_unsigned(9081,N);
          when 642 =>   sin_data_int <= to_unsigned(13650,N); cos_data_int <= to_unsigned(9060,N);
          when 643 =>   sin_data_int <= to_unsigned(13664,N); cos_data_int <= to_unsigned(9039,N);
          when 644 =>   sin_data_int <= to_unsigned(13678,N); cos_data_int <= to_unsigned(9018,N);
          when 645 =>   sin_data_int <= to_unsigned(13692,N); cos_data_int <= to_unsigned(8997,N);
          when 646 =>   sin_data_int <= to_unsigned(13705,N); cos_data_int <= to_unsigned(8976,N);
          when 647 =>   sin_data_int <= to_unsigned(13719,N); cos_data_int <= to_unsigned(8955,N);
          when 648 =>   sin_data_int <= to_unsigned(13733,N); cos_data_int <= to_unsigned(8934,N);
          when 649 =>   sin_data_int <= to_unsigned(13747,N); cos_data_int <= to_unsigned(8913,N);
          when 650 =>   sin_data_int <= to_unsigned(13760,N); cos_data_int <= to_unsigned(8892,N);
          when 651 =>   sin_data_int <= to_unsigned(13774,N); cos_data_int <= to_unsigned(8871,N);
          when 652 =>   sin_data_int <= to_unsigned(13788,N); cos_data_int <= to_unsigned(8850,N);
          when 653 =>   sin_data_int <= to_unsigned(13801,N); cos_data_int <= to_unsigned(8829,N);
          when 654 =>   sin_data_int <= to_unsigned(13815,N); cos_data_int <= to_unsigned(8807,N);
          when 655 =>   sin_data_int <= to_unsigned(13828,N); cos_data_int <= to_unsigned(8786,N);
          when 656 =>   sin_data_int <= to_unsigned(13842,N); cos_data_int <= to_unsigned(8765,N);
          when 657 =>   sin_data_int <= to_unsigned(13855,N); cos_data_int <= to_unsigned(8744,N);
          when 658 =>   sin_data_int <= to_unsigned(13868,N); cos_data_int <= to_unsigned(8722,N);
          when 659 =>   sin_data_int <= to_unsigned(13882,N); cos_data_int <= to_unsigned(8701,N);
          when 660 =>   sin_data_int <= to_unsigned(13895,N); cos_data_int <= to_unsigned(8680,N);
          when 661 =>   sin_data_int <= to_unsigned(13908,N); cos_data_int <= to_unsigned(8658,N);
          when 662 =>   sin_data_int <= to_unsigned(13922,N); cos_data_int <= to_unsigned(8637,N);
          when 663 =>   sin_data_int <= to_unsigned(13935,N); cos_data_int <= to_unsigned(8616,N);
          when 664 =>   sin_data_int <= to_unsigned(13948,N); cos_data_int <= to_unsigned(8594,N);
          when 665 =>   sin_data_int <= to_unsigned(13961,N); cos_data_int <= to_unsigned(8573,N);
          when 666 =>   sin_data_int <= to_unsigned(13974,N); cos_data_int <= to_unsigned(8552,N);
          when 667 =>   sin_data_int <= to_unsigned(13988,N); cos_data_int <= to_unsigned(8530,N);
          when 668 =>   sin_data_int <= to_unsigned(14001,N); cos_data_int <= to_unsigned(8509,N);
          when 669 =>   sin_data_int <= to_unsigned(14014,N); cos_data_int <= to_unsigned(8487,N);
          when 670 =>   sin_data_int <= to_unsigned(14027,N); cos_data_int <= to_unsigned(8466,N);
          when 671 =>   sin_data_int <= to_unsigned(14040,N); cos_data_int <= to_unsigned(8444,N);
          when 672 =>   sin_data_int <= to_unsigned(14053,N); cos_data_int <= to_unsigned(8423,N);
          when 673 =>   sin_data_int <= to_unsigned(14065,N); cos_data_int <= to_unsigned(8401,N);
          when 674 =>   sin_data_int <= to_unsigned(14078,N); cos_data_int <= to_unsigned(8379,N);
          when 675 =>   sin_data_int <= to_unsigned(14091,N); cos_data_int <= to_unsigned(8358,N);
          when 676 =>   sin_data_int <= to_unsigned(14104,N); cos_data_int <= to_unsigned(8336,N);
          when 677 =>   sin_data_int <= to_unsigned(14117,N); cos_data_int <= to_unsigned(8315,N);
          when 678 =>   sin_data_int <= to_unsigned(14129,N); cos_data_int <= to_unsigned(8293,N);
          when 679 =>   sin_data_int <= to_unsigned(14142,N); cos_data_int <= to_unsigned(8271,N);
          when 680 =>   sin_data_int <= to_unsigned(14155,N); cos_data_int <= to_unsigned(8249,N);
          when 681 =>   sin_data_int <= to_unsigned(14167,N); cos_data_int <= to_unsigned(8228,N);
          when 682 =>   sin_data_int <= to_unsigned(14180,N); cos_data_int <= to_unsigned(8206,N);
          when 683 =>   sin_data_int <= to_unsigned(14193,N); cos_data_int <= to_unsigned(8184,N);
          when 684 =>   sin_data_int <= to_unsigned(14205,N); cos_data_int <= to_unsigned(8162,N);
          when 685 =>   sin_data_int <= to_unsigned(14218,N); cos_data_int <= to_unsigned(8141,N);
          when 686 =>   sin_data_int <= to_unsigned(14230,N); cos_data_int <= to_unsigned(8119,N);
          when 687 =>   sin_data_int <= to_unsigned(14243,N); cos_data_int <= to_unsigned(8097,N);
          when 688 =>   sin_data_int <= to_unsigned(14255,N); cos_data_int <= to_unsigned(8075,N);
          when 689 =>   sin_data_int <= to_unsigned(14267,N); cos_data_int <= to_unsigned(8053,N);
          when 690 =>   sin_data_int <= to_unsigned(14280,N); cos_data_int <= to_unsigned(8031,N);
          when 691 =>   sin_data_int <= to_unsigned(14292,N); cos_data_int <= to_unsigned(8009,N);
          when 692 =>   sin_data_int <= to_unsigned(14304,N); cos_data_int <= to_unsigned(7988,N);
          when 693 =>   sin_data_int <= to_unsigned(14317,N); cos_data_int <= to_unsigned(7966,N);
          when 694 =>   sin_data_int <= to_unsigned(14329,N); cos_data_int <= to_unsigned(7944,N);
          when 695 =>   sin_data_int <= to_unsigned(14341,N); cos_data_int <= to_unsigned(7922,N);
          when 696 =>   sin_data_int <= to_unsigned(14353,N); cos_data_int <= to_unsigned(7900,N);
          when 697 =>   sin_data_int <= to_unsigned(14365,N); cos_data_int <= to_unsigned(7878,N);
          when 698 =>   sin_data_int <= to_unsigned(14377,N); cos_data_int <= to_unsigned(7856,N);
          when 699 =>   sin_data_int <= to_unsigned(14389,N); cos_data_int <= to_unsigned(7833,N);
          when 700 =>   sin_data_int <= to_unsigned(14401,N); cos_data_int <= to_unsigned(7811,N);
          when 701 =>   sin_data_int <= to_unsigned(14413,N); cos_data_int <= to_unsigned(7789,N);
          when 702 =>   sin_data_int <= to_unsigned(14425,N); cos_data_int <= to_unsigned(7767,N);
          when 703 =>   sin_data_int <= to_unsigned(14437,N); cos_data_int <= to_unsigned(7745,N);
          when 704 =>   sin_data_int <= to_unsigned(14449,N); cos_data_int <= to_unsigned(7723,N);
          when 705 =>   sin_data_int <= to_unsigned(14461,N); cos_data_int <= to_unsigned(7701,N);
          when 706 =>   sin_data_int <= to_unsigned(14473,N); cos_data_int <= to_unsigned(7678,N);
          when 707 =>   sin_data_int <= to_unsigned(14484,N); cos_data_int <= to_unsigned(7656,N);
          when 708 =>   sin_data_int <= to_unsigned(14496,N); cos_data_int <= to_unsigned(7634,N);
          when 709 =>   sin_data_int <= to_unsigned(14508,N); cos_data_int <= to_unsigned(7612,N);
          when 710 =>   sin_data_int <= to_unsigned(14519,N); cos_data_int <= to_unsigned(7590,N);
          when 711 =>   sin_data_int <= to_unsigned(14531,N); cos_data_int <= to_unsigned(7567,N);
          when 712 =>   sin_data_int <= to_unsigned(14543,N); cos_data_int <= to_unsigned(7545,N);
          when 713 =>   sin_data_int <= to_unsigned(14554,N); cos_data_int <= to_unsigned(7523,N);
          when 714 =>   sin_data_int <= to_unsigned(14566,N); cos_data_int <= to_unsigned(7500,N);
          when 715 =>   sin_data_int <= to_unsigned(14577,N); cos_data_int <= to_unsigned(7478,N);
          when 716 =>   sin_data_int <= to_unsigned(14589,N); cos_data_int <= to_unsigned(7456,N);
          when 717 =>   sin_data_int <= to_unsigned(14600,N); cos_data_int <= to_unsigned(7433,N);
          when 718 =>   sin_data_int <= to_unsigned(14611,N); cos_data_int <= to_unsigned(7411,N);
          when 719 =>   sin_data_int <= to_unsigned(14623,N); cos_data_int <= to_unsigned(7388,N);
          when 720 =>   sin_data_int <= to_unsigned(14634,N); cos_data_int <= to_unsigned(7366,N);
          when 721 =>   sin_data_int <= to_unsigned(14645,N); cos_data_int <= to_unsigned(7343,N);
          when 722 =>   sin_data_int <= to_unsigned(14657,N); cos_data_int <= to_unsigned(7321,N);
          when 723 =>   sin_data_int <= to_unsigned(14668,N); cos_data_int <= to_unsigned(7299,N);
          when 724 =>   sin_data_int <= to_unsigned(14679,N); cos_data_int <= to_unsigned(7276,N);
          when 725 =>   sin_data_int <= to_unsigned(14690,N); cos_data_int <= to_unsigned(7253,N);
          when 726 =>   sin_data_int <= to_unsigned(14701,N); cos_data_int <= to_unsigned(7231,N);
          when 727 =>   sin_data_int <= to_unsigned(14712,N); cos_data_int <= to_unsigned(7208,N);
          when 728 =>   sin_data_int <= to_unsigned(14723,N); cos_data_int <= to_unsigned(7186,N);
          when 729 =>   sin_data_int <= to_unsigned(14734,N); cos_data_int <= to_unsigned(7163,N);
          when 730 =>   sin_data_int <= to_unsigned(14745,N); cos_data_int <= to_unsigned(7141,N);
          when 731 =>   sin_data_int <= to_unsigned(14756,N); cos_data_int <= to_unsigned(7118,N);
          when 732 =>   sin_data_int <= to_unsigned(14767,N); cos_data_int <= to_unsigned(7095,N);
          when 733 =>   sin_data_int <= to_unsigned(14778,N); cos_data_int <= to_unsigned(7073,N);
          when 734 =>   sin_data_int <= to_unsigned(14789,N); cos_data_int <= to_unsigned(7050,N);
          when 735 =>   sin_data_int <= to_unsigned(14800,N); cos_data_int <= to_unsigned(7027,N);
          when 736 =>   sin_data_int <= to_unsigned(14810,N); cos_data_int <= to_unsigned(7005,N);
          when 737 =>   sin_data_int <= to_unsigned(14821,N); cos_data_int <= to_unsigned(6982,N);
          when 738 =>   sin_data_int <= to_unsigned(14832,N); cos_data_int <= to_unsigned(6959,N);
          when 739 =>   sin_data_int <= to_unsigned(14843,N); cos_data_int <= to_unsigned(6936,N);
          when 740 =>   sin_data_int <= to_unsigned(14853,N); cos_data_int <= to_unsigned(6914,N);
          when 741 =>   sin_data_int <= to_unsigned(14864,N); cos_data_int <= to_unsigned(6891,N);
          when 742 =>   sin_data_int <= to_unsigned(14874,N); cos_data_int <= to_unsigned(6868,N);
          when 743 =>   sin_data_int <= to_unsigned(14885,N); cos_data_int <= to_unsigned(6845,N);
          when 744 =>   sin_data_int <= to_unsigned(14895,N); cos_data_int <= to_unsigned(6822,N);
          when 745 =>   sin_data_int <= to_unsigned(14906,N); cos_data_int <= to_unsigned(6799,N);
          when 746 =>   sin_data_int <= to_unsigned(14916,N); cos_data_int <= to_unsigned(6777,N);
          when 747 =>   sin_data_int <= to_unsigned(14927,N); cos_data_int <= to_unsigned(6754,N);
          when 748 =>   sin_data_int <= to_unsigned(14937,N); cos_data_int <= to_unsigned(6731,N);
          when 749 =>   sin_data_int <= to_unsigned(14947,N); cos_data_int <= to_unsigned(6708,N);
          when 750 =>   sin_data_int <= to_unsigned(14957,N); cos_data_int <= to_unsigned(6685,N);
          when 751 =>   sin_data_int <= to_unsigned(14968,N); cos_data_int <= to_unsigned(6662,N);
          when 752 =>   sin_data_int <= to_unsigned(14978,N); cos_data_int <= to_unsigned(6639,N);
          when 753 =>   sin_data_int <= to_unsigned(14988,N); cos_data_int <= to_unsigned(6616,N);
          when 754 =>   sin_data_int <= to_unsigned(14998,N); cos_data_int <= to_unsigned(6593,N);
          when 755 =>   sin_data_int <= to_unsigned(15008,N); cos_data_int <= to_unsigned(6570,N);
          when 756 =>   sin_data_int <= to_unsigned(15018,N); cos_data_int <= to_unsigned(6547,N);
          when 757 =>   sin_data_int <= to_unsigned(15028,N); cos_data_int <= to_unsigned(6524,N);
          when 758 =>   sin_data_int <= to_unsigned(15038,N); cos_data_int <= to_unsigned(6501,N);
          when 759 =>   sin_data_int <= to_unsigned(15048,N); cos_data_int <= to_unsigned(6478,N);
          when 760 =>   sin_data_int <= to_unsigned(15058,N); cos_data_int <= to_unsigned(6455,N);
          when 761 =>   sin_data_int <= to_unsigned(15068,N); cos_data_int <= to_unsigned(6432,N);
          when 762 =>   sin_data_int <= to_unsigned(15078,N); cos_data_int <= to_unsigned(6408,N);
          when 763 =>   sin_data_int <= to_unsigned(15088,N); cos_data_int <= to_unsigned(6385,N);
          when 764 =>   sin_data_int <= to_unsigned(15098,N); cos_data_int <= to_unsigned(6362,N);
          when 765 =>   sin_data_int <= to_unsigned(15107,N); cos_data_int <= to_unsigned(6339,N);
          when 766 =>   sin_data_int <= to_unsigned(15117,N); cos_data_int <= to_unsigned(6316,N);
          when 767 =>   sin_data_int <= to_unsigned(15127,N); cos_data_int <= to_unsigned(6293,N);
          when 768 =>   sin_data_int <= to_unsigned(15136,N); cos_data_int <= to_unsigned(6269,N);
          when 769 =>   sin_data_int <= to_unsigned(15146,N); cos_data_int <= to_unsigned(6246,N);
          when 770 =>   sin_data_int <= to_unsigned(15156,N); cos_data_int <= to_unsigned(6223,N);
          when 771 =>   sin_data_int <= to_unsigned(15165,N); cos_data_int <= to_unsigned(6200,N);
          when 772 =>   sin_data_int <= to_unsigned(15175,N); cos_data_int <= to_unsigned(6176,N);
          when 773 =>   sin_data_int <= to_unsigned(15184,N); cos_data_int <= to_unsigned(6153,N);
          when 774 =>   sin_data_int <= to_unsigned(15193,N); cos_data_int <= to_unsigned(6130,N);
          when 775 =>   sin_data_int <= to_unsigned(15203,N); cos_data_int <= to_unsigned(6106,N);
          when 776 =>   sin_data_int <= to_unsigned(15212,N); cos_data_int <= to_unsigned(6083,N);
          when 777 =>   sin_data_int <= to_unsigned(15221,N); cos_data_int <= to_unsigned(6060,N);
          when 778 =>   sin_data_int <= to_unsigned(15231,N); cos_data_int <= to_unsigned(6036,N);
          when 779 =>   sin_data_int <= to_unsigned(15240,N); cos_data_int <= to_unsigned(6013,N);
          when 780 =>   sin_data_int <= to_unsigned(15249,N); cos_data_int <= to_unsigned(5990,N);
          when 781 =>   sin_data_int <= to_unsigned(15258,N); cos_data_int <= to_unsigned(5966,N);
          when 782 =>   sin_data_int <= to_unsigned(15267,N); cos_data_int <= to_unsigned(5943,N);
          when 783 =>   sin_data_int <= to_unsigned(15277,N); cos_data_int <= to_unsigned(5919,N);
          when 784 =>   sin_data_int <= to_unsigned(15286,N); cos_data_int <= to_unsigned(5896,N);
          when 785 =>   sin_data_int <= to_unsigned(15295,N); cos_data_int <= to_unsigned(5873,N);
          when 786 =>   sin_data_int <= to_unsigned(15304,N); cos_data_int <= to_unsigned(5849,N);
          when 787 =>   sin_data_int <= to_unsigned(15313,N); cos_data_int <= to_unsigned(5826,N);
          when 788 =>   sin_data_int <= to_unsigned(15322,N); cos_data_int <= to_unsigned(5802,N);
          when 789 =>   sin_data_int <= to_unsigned(15330,N); cos_data_int <= to_unsigned(5779,N);
          when 790 =>   sin_data_int <= to_unsigned(15339,N); cos_data_int <= to_unsigned(5755,N);
          when 791 =>   sin_data_int <= to_unsigned(15348,N); cos_data_int <= to_unsigned(5732,N);
          when 792 =>   sin_data_int <= to_unsigned(15357,N); cos_data_int <= to_unsigned(5708,N);
          when 793 =>   sin_data_int <= to_unsigned(15366,N); cos_data_int <= to_unsigned(5684,N);
          when 794 =>   sin_data_int <= to_unsigned(15374,N); cos_data_int <= to_unsigned(5661,N);
          when 795 =>   sin_data_int <= to_unsigned(15383,N); cos_data_int <= to_unsigned(5637,N);
          when 796 =>   sin_data_int <= to_unsigned(15392,N); cos_data_int <= to_unsigned(5614,N);
          when 797 =>   sin_data_int <= to_unsigned(15400,N); cos_data_int <= to_unsigned(5590,N);
          when 798 =>   sin_data_int <= to_unsigned(15409,N); cos_data_int <= to_unsigned(5566,N);
          when 799 =>   sin_data_int <= to_unsigned(15417,N); cos_data_int <= to_unsigned(5543,N);
          when 800 =>   sin_data_int <= to_unsigned(15426,N); cos_data_int <= to_unsigned(5519,N);
          when 801 =>   sin_data_int <= to_unsigned(15434,N); cos_data_int <= to_unsigned(5495,N);
          when 802 =>   sin_data_int <= to_unsigned(15443,N); cos_data_int <= to_unsigned(5472,N);
          when 803 =>   sin_data_int <= to_unsigned(15451,N); cos_data_int <= to_unsigned(5448,N);
          when 804 =>   sin_data_int <= to_unsigned(15459,N); cos_data_int <= to_unsigned(5424,N);
          when 805 =>   sin_data_int <= to_unsigned(15468,N); cos_data_int <= to_unsigned(5401,N);
          when 806 =>   sin_data_int <= to_unsigned(15476,N); cos_data_int <= to_unsigned(5377,N);
          when 807 =>   sin_data_int <= to_unsigned(15484,N); cos_data_int <= to_unsigned(5353,N);
          when 808 =>   sin_data_int <= to_unsigned(15492,N); cos_data_int <= to_unsigned(5329,N);
          when 809 =>   sin_data_int <= to_unsigned(15500,N); cos_data_int <= to_unsigned(5306,N);
          when 810 =>   sin_data_int <= to_unsigned(15509,N); cos_data_int <= to_unsigned(5282,N);
          when 811 =>   sin_data_int <= to_unsigned(15517,N); cos_data_int <= to_unsigned(5258,N);
          when 812 =>   sin_data_int <= to_unsigned(15525,N); cos_data_int <= to_unsigned(5234,N);
          when 813 =>   sin_data_int <= to_unsigned(15533,N); cos_data_int <= to_unsigned(5210,N);
          when 814 =>   sin_data_int <= to_unsigned(15541,N); cos_data_int <= to_unsigned(5187,N);
          when 815 =>   sin_data_int <= to_unsigned(15549,N); cos_data_int <= to_unsigned(5163,N);
          when 816 =>   sin_data_int <= to_unsigned(15557,N); cos_data_int <= to_unsigned(5139,N);
          when 817 =>   sin_data_int <= to_unsigned(15564,N); cos_data_int <= to_unsigned(5115,N);
          when 818 =>   sin_data_int <= to_unsigned(15572,N); cos_data_int <= to_unsigned(5091,N);
          when 819 =>   sin_data_int <= to_unsigned(15580,N); cos_data_int <= to_unsigned(5067,N);
          when 820 =>   sin_data_int <= to_unsigned(15588,N); cos_data_int <= to_unsigned(5043,N);
          when 821 =>   sin_data_int <= to_unsigned(15596,N); cos_data_int <= to_unsigned(5019,N);
          when 822 =>   sin_data_int <= to_unsigned(15603,N); cos_data_int <= to_unsigned(4995,N);
          when 823 =>   sin_data_int <= to_unsigned(15611,N); cos_data_int <= to_unsigned(4972,N);
          when 824 =>   sin_data_int <= to_unsigned(15618,N); cos_data_int <= to_unsigned(4948,N);
          when 825 =>   sin_data_int <= to_unsigned(15626,N); cos_data_int <= to_unsigned(4924,N);
          when 826 =>   sin_data_int <= to_unsigned(15634,N); cos_data_int <= to_unsigned(4900,N);
          when 827 =>   sin_data_int <= to_unsigned(15641,N); cos_data_int <= to_unsigned(4876,N);
          when 828 =>   sin_data_int <= to_unsigned(15649,N); cos_data_int <= to_unsigned(4852,N);
          when 829 =>   sin_data_int <= to_unsigned(15656,N); cos_data_int <= to_unsigned(4828,N);
          when 830 =>   sin_data_int <= to_unsigned(15663,N); cos_data_int <= to_unsigned(4804,N);
          when 831 =>   sin_data_int <= to_unsigned(15671,N); cos_data_int <= to_unsigned(4780,N);
          when 832 =>   sin_data_int <= to_unsigned(15678,N); cos_data_int <= to_unsigned(4756,N);
          when 833 =>   sin_data_int <= to_unsigned(15685,N); cos_data_int <= to_unsigned(4731,N);
          when 834 =>   sin_data_int <= to_unsigned(15693,N); cos_data_int <= to_unsigned(4707,N);
          when 835 =>   sin_data_int <= to_unsigned(15700,N); cos_data_int <= to_unsigned(4683,N);
          when 836 =>   sin_data_int <= to_unsigned(15707,N); cos_data_int <= to_unsigned(4659,N);
          when 837 =>   sin_data_int <= to_unsigned(15714,N); cos_data_int <= to_unsigned(4635,N);
          when 838 =>   sin_data_int <= to_unsigned(15721,N); cos_data_int <= to_unsigned(4611,N);
          when 839 =>   sin_data_int <= to_unsigned(15728,N); cos_data_int <= to_unsigned(4587,N);
          when 840 =>   sin_data_int <= to_unsigned(15735,N); cos_data_int <= to_unsigned(4563,N);
          when 841 =>   sin_data_int <= to_unsigned(15742,N); cos_data_int <= to_unsigned(4539,N);
          when 842 =>   sin_data_int <= to_unsigned(15749,N); cos_data_int <= to_unsigned(4514,N);
          when 843 =>   sin_data_int <= to_unsigned(15756,N); cos_data_int <= to_unsigned(4490,N);
          when 844 =>   sin_data_int <= to_unsigned(15763,N); cos_data_int <= to_unsigned(4466,N);
          when 845 =>   sin_data_int <= to_unsigned(15770,N); cos_data_int <= to_unsigned(4442,N);
          when 846 =>   sin_data_int <= to_unsigned(15777,N); cos_data_int <= to_unsigned(4418,N);
          when 847 =>   sin_data_int <= to_unsigned(15783,N); cos_data_int <= to_unsigned(4394,N);
          when 848 =>   sin_data_int <= to_unsigned(15790,N); cos_data_int <= to_unsigned(4369,N);
          when 849 =>   sin_data_int <= to_unsigned(15797,N); cos_data_int <= to_unsigned(4345,N);
          when 850 =>   sin_data_int <= to_unsigned(15803,N); cos_data_int <= to_unsigned(4321,N);
          when 851 =>   sin_data_int <= to_unsigned(15810,N); cos_data_int <= to_unsigned(4297,N);
          when 852 =>   sin_data_int <= to_unsigned(15817,N); cos_data_int <= to_unsigned(4272,N);
          when 853 =>   sin_data_int <= to_unsigned(15823,N); cos_data_int <= to_unsigned(4248,N);
          when 854 =>   sin_data_int <= to_unsigned(15830,N); cos_data_int <= to_unsigned(4224,N);
          when 855 =>   sin_data_int <= to_unsigned(15836,N); cos_data_int <= to_unsigned(4200,N);
          when 856 =>   sin_data_int <= to_unsigned(15842,N); cos_data_int <= to_unsigned(4175,N);
          when 857 =>   sin_data_int <= to_unsigned(15849,N); cos_data_int <= to_unsigned(4151,N);
          when 858 =>   sin_data_int <= to_unsigned(15855,N); cos_data_int <= to_unsigned(4127,N);
          when 859 =>   sin_data_int <= to_unsigned(15861,N); cos_data_int <= to_unsigned(4102,N);
          when 860 =>   sin_data_int <= to_unsigned(15868,N); cos_data_int <= to_unsigned(4078,N);
          when 861 =>   sin_data_int <= to_unsigned(15874,N); cos_data_int <= to_unsigned(4054,N);
          when 862 =>   sin_data_int <= to_unsigned(15880,N); cos_data_int <= to_unsigned(4029,N);
          when 863 =>   sin_data_int <= to_unsigned(15886,N); cos_data_int <= to_unsigned(4005,N);
          when 864 =>   sin_data_int <= to_unsigned(15892,N); cos_data_int <= to_unsigned(3980,N);
          when 865 =>   sin_data_int <= to_unsigned(15899,N); cos_data_int <= to_unsigned(3956,N);
          when 866 =>   sin_data_int <= to_unsigned(15905,N); cos_data_int <= to_unsigned(3932,N);
          when 867 =>   sin_data_int <= to_unsigned(15911,N); cos_data_int <= to_unsigned(3907,N);
          when 868 =>   sin_data_int <= to_unsigned(15917,N); cos_data_int <= to_unsigned(3883,N);
          when 869 =>   sin_data_int <= to_unsigned(15923,N); cos_data_int <= to_unsigned(3858,N);
          when 870 =>   sin_data_int <= to_unsigned(15928,N); cos_data_int <= to_unsigned(3834,N);
          when 871 =>   sin_data_int <= to_unsigned(15934,N); cos_data_int <= to_unsigned(3810,N);
          when 872 =>   sin_data_int <= to_unsigned(15940,N); cos_data_int <= to_unsigned(3785,N);
          when 873 =>   sin_data_int <= to_unsigned(15946,N); cos_data_int <= to_unsigned(3761,N);
          when 874 =>   sin_data_int <= to_unsigned(15952,N); cos_data_int <= to_unsigned(3736,N);
          when 875 =>   sin_data_int <= to_unsigned(15957,N); cos_data_int <= to_unsigned(3712,N);
          when 876 =>   sin_data_int <= to_unsigned(15963,N); cos_data_int <= to_unsigned(3687,N);
          when 877 =>   sin_data_int <= to_unsigned(15969,N); cos_data_int <= to_unsigned(3663,N);
          when 878 =>   sin_data_int <= to_unsigned(15974,N); cos_data_int <= to_unsigned(3638,N);
          when 879 =>   sin_data_int <= to_unsigned(15980,N); cos_data_int <= to_unsigned(3614,N);
          when 880 =>   sin_data_int <= to_unsigned(15985,N); cos_data_int <= to_unsigned(3589,N);
          when 881 =>   sin_data_int <= to_unsigned(15991,N); cos_data_int <= to_unsigned(3565,N);
          when 882 =>   sin_data_int <= to_unsigned(15996,N); cos_data_int <= to_unsigned(3540,N);
          when 883 =>   sin_data_int <= to_unsigned(16002,N); cos_data_int <= to_unsigned(3516,N);
          when 884 =>   sin_data_int <= to_unsigned(16007,N); cos_data_int <= to_unsigned(3491,N);
          when 885 =>   sin_data_int <= to_unsigned(16012,N); cos_data_int <= to_unsigned(3467,N);
          when 886 =>   sin_data_int <= to_unsigned(16018,N); cos_data_int <= to_unsigned(3442,N);
          when 887 =>   sin_data_int <= to_unsigned(16023,N); cos_data_int <= to_unsigned(3417,N);
          when 888 =>   sin_data_int <= to_unsigned(16028,N); cos_data_int <= to_unsigned(3393,N);
          when 889 =>   sin_data_int <= to_unsigned(16033,N); cos_data_int <= to_unsigned(3368,N);
          when 890 =>   sin_data_int <= to_unsigned(16039,N); cos_data_int <= to_unsigned(3344,N);
          when 891 =>   sin_data_int <= to_unsigned(16044,N); cos_data_int <= to_unsigned(3319,N);
          when 892 =>   sin_data_int <= to_unsigned(16049,N); cos_data_int <= to_unsigned(3294,N);
          when 893 =>   sin_data_int <= to_unsigned(16054,N); cos_data_int <= to_unsigned(3270,N);
          when 894 =>   sin_data_int <= to_unsigned(16059,N); cos_data_int <= to_unsigned(3245,N);
          when 895 =>   sin_data_int <= to_unsigned(16064,N); cos_data_int <= to_unsigned(3221,N);
          when 896 =>   sin_data_int <= to_unsigned(16069,N); cos_data_int <= to_unsigned(3196,N);
          when 897 =>   sin_data_int <= to_unsigned(16074,N); cos_data_int <= to_unsigned(3171,N);
          when 898 =>   sin_data_int <= to_unsigned(16078,N); cos_data_int <= to_unsigned(3147,N);
          when 899 =>   sin_data_int <= to_unsigned(16083,N); cos_data_int <= to_unsigned(3122,N);
          when 900 =>   sin_data_int <= to_unsigned(16088,N); cos_data_int <= to_unsigned(3097,N);
          when 901 =>   sin_data_int <= to_unsigned(16093,N); cos_data_int <= to_unsigned(3073,N);
          when 902 =>   sin_data_int <= to_unsigned(16097,N); cos_data_int <= to_unsigned(3048,N);
          when 903 =>   sin_data_int <= to_unsigned(16102,N); cos_data_int <= to_unsigned(3023,N);
          when 904 =>   sin_data_int <= to_unsigned(16107,N); cos_data_int <= to_unsigned(2998,N);
          when 905 =>   sin_data_int <= to_unsigned(16111,N); cos_data_int <= to_unsigned(2974,N);
          when 906 =>   sin_data_int <= to_unsigned(16116,N); cos_data_int <= to_unsigned(2949,N);
          when 907 =>   sin_data_int <= to_unsigned(16120,N); cos_data_int <= to_unsigned(2924,N);
          when 908 =>   sin_data_int <= to_unsigned(16125,N); cos_data_int <= to_unsigned(2900,N);
          when 909 =>   sin_data_int <= to_unsigned(16129,N); cos_data_int <= to_unsigned(2875,N);
          when 910 =>   sin_data_int <= to_unsigned(16134,N); cos_data_int <= to_unsigned(2850,N);
          when 911 =>   sin_data_int <= to_unsigned(16138,N); cos_data_int <= to_unsigned(2825,N);
          when 912 =>   sin_data_int <= to_unsigned(16142,N); cos_data_int <= to_unsigned(2801,N);
          when 913 =>   sin_data_int <= to_unsigned(16147,N); cos_data_int <= to_unsigned(2776,N);
          when 914 =>   sin_data_int <= to_unsigned(16151,N); cos_data_int <= to_unsigned(2751,N);
          when 915 =>   sin_data_int <= to_unsigned(16155,N); cos_data_int <= to_unsigned(2726,N);
          when 916 =>   sin_data_int <= to_unsigned(16159,N); cos_data_int <= to_unsigned(2701,N);
          when 917 =>   sin_data_int <= to_unsigned(16163,N); cos_data_int <= to_unsigned(2677,N);
          when 918 =>   sin_data_int <= to_unsigned(16167,N); cos_data_int <= to_unsigned(2652,N);
          when 919 =>   sin_data_int <= to_unsigned(16171,N); cos_data_int <= to_unsigned(2627,N);
          when 920 =>   sin_data_int <= to_unsigned(16175,N); cos_data_int <= to_unsigned(2602,N);
          when 921 =>   sin_data_int <= to_unsigned(16179,N); cos_data_int <= to_unsigned(2577,N);
          when 922 =>   sin_data_int <= to_unsigned(16183,N); cos_data_int <= to_unsigned(2553,N);
          when 923 =>   sin_data_int <= to_unsigned(16187,N); cos_data_int <= to_unsigned(2528,N);
          when 924 =>   sin_data_int <= to_unsigned(16191,N); cos_data_int <= to_unsigned(2503,N);
          when 925 =>   sin_data_int <= to_unsigned(16195,N); cos_data_int <= to_unsigned(2478,N);
          when 926 =>   sin_data_int <= to_unsigned(16199,N); cos_data_int <= to_unsigned(2453,N);
          when 927 =>   sin_data_int <= to_unsigned(16202,N); cos_data_int <= to_unsigned(2428,N);
          when 928 =>   sin_data_int <= to_unsigned(16206,N); cos_data_int <= to_unsigned(2404,N);
          when 929 =>   sin_data_int <= to_unsigned(16210,N); cos_data_int <= to_unsigned(2379,N);
          when 930 =>   sin_data_int <= to_unsigned(16213,N); cos_data_int <= to_unsigned(2354,N);
          when 931 =>   sin_data_int <= to_unsigned(16217,N); cos_data_int <= to_unsigned(2329,N);
          when 932 =>   sin_data_int <= to_unsigned(16221,N); cos_data_int <= to_unsigned(2304,N);
          when 933 =>   sin_data_int <= to_unsigned(16224,N); cos_data_int <= to_unsigned(2279,N);
          when 934 =>   sin_data_int <= to_unsigned(16228,N); cos_data_int <= to_unsigned(2254,N);
          when 935 =>   sin_data_int <= to_unsigned(16231,N); cos_data_int <= to_unsigned(2229,N);
          when 936 =>   sin_data_int <= to_unsigned(16234,N); cos_data_int <= to_unsigned(2204,N);
          when 937 =>   sin_data_int <= to_unsigned(16238,N); cos_data_int <= to_unsigned(2180,N);
          when 938 =>   sin_data_int <= to_unsigned(16241,N); cos_data_int <= to_unsigned(2155,N);
          when 939 =>   sin_data_int <= to_unsigned(16244,N); cos_data_int <= to_unsigned(2130,N);
          when 940 =>   sin_data_int <= to_unsigned(16248,N); cos_data_int <= to_unsigned(2105,N);
          when 941 =>   sin_data_int <= to_unsigned(16251,N); cos_data_int <= to_unsigned(2080,N);
          when 942 =>   sin_data_int <= to_unsigned(16254,N); cos_data_int <= to_unsigned(2055,N);
          when 943 =>   sin_data_int <= to_unsigned(16257,N); cos_data_int <= to_unsigned(2030,N);
          when 944 =>   sin_data_int <= to_unsigned(16260,N); cos_data_int <= to_unsigned(2005,N);
          when 945 =>   sin_data_int <= to_unsigned(16263,N); cos_data_int <= to_unsigned(1980,N);
          when 946 =>   sin_data_int <= to_unsigned(16266,N); cos_data_int <= to_unsigned(1955,N);
          when 947 =>   sin_data_int <= to_unsigned(16269,N); cos_data_int <= to_unsigned(1930,N);
          when 948 =>   sin_data_int <= to_unsigned(16272,N); cos_data_int <= to_unsigned(1905,N);
          when 949 =>   sin_data_int <= to_unsigned(16275,N); cos_data_int <= to_unsigned(1880,N);
          when 950 =>   sin_data_int <= to_unsigned(16278,N); cos_data_int <= to_unsigned(1855,N);
          when 951 =>   sin_data_int <= to_unsigned(16281,N); cos_data_int <= to_unsigned(1830,N);
          when 952 =>   sin_data_int <= to_unsigned(16284,N); cos_data_int <= to_unsigned(1805,N);
          when 953 =>   sin_data_int <= to_unsigned(16286,N); cos_data_int <= to_unsigned(1780,N);
          when 954 =>   sin_data_int <= to_unsigned(16289,N); cos_data_int <= to_unsigned(1755,N);
          when 955 =>   sin_data_int <= to_unsigned(16292,N); cos_data_int <= to_unsigned(1730,N);
          when 956 =>   sin_data_int <= to_unsigned(16294,N); cos_data_int <= to_unsigned(1705,N);
          when 957 =>   sin_data_int <= to_unsigned(16297,N); cos_data_int <= to_unsigned(1680,N);
          when 958 =>   sin_data_int <= to_unsigned(16300,N); cos_data_int <= to_unsigned(1655,N);
          when 959 =>   sin_data_int <= to_unsigned(16302,N); cos_data_int <= to_unsigned(1630,N);
          when 960 =>   sin_data_int <= to_unsigned(16305,N); cos_data_int <= to_unsigned(1605,N);
          when 961 =>   sin_data_int <= to_unsigned(16307,N); cos_data_int <= to_unsigned(1580,N);
          when 962 =>   sin_data_int <= to_unsigned(16309,N); cos_data_int <= to_unsigned(1555,N);
          when 963 =>   sin_data_int <= to_unsigned(16312,N); cos_data_int <= to_unsigned(1530,N);
          when 964 =>   sin_data_int <= to_unsigned(16314,N); cos_data_int <= to_unsigned(1505,N);
          when 965 =>   sin_data_int <= to_unsigned(16316,N); cos_data_int <= to_unsigned(1480,N);
          when 966 =>   sin_data_int <= to_unsigned(16319,N); cos_data_int <= to_unsigned(1455,N);
          when 967 =>   sin_data_int <= to_unsigned(16321,N); cos_data_int <= to_unsigned(1430,N);
          when 968 =>   sin_data_int <= to_unsigned(16323,N); cos_data_int <= to_unsigned(1405,N);
          when 969 =>   sin_data_int <= to_unsigned(16325,N); cos_data_int <= to_unsigned(1380,N);
          when 970 =>   sin_data_int <= to_unsigned(16327,N); cos_data_int <= to_unsigned(1355,N);
          when 971 =>   sin_data_int <= to_unsigned(16329,N); cos_data_int <= to_unsigned(1330,N);
          when 972 =>   sin_data_int <= to_unsigned(16331,N); cos_data_int <= to_unsigned(1305,N);
          when 973 =>   sin_data_int <= to_unsigned(16333,N); cos_data_int <= to_unsigned(1280,N);
          when 974 =>   sin_data_int <= to_unsigned(16335,N); cos_data_int <= to_unsigned(1255,N);
          when 975 =>   sin_data_int <= to_unsigned(16337,N); cos_data_int <= to_unsigned(1230,N);
          when 976 =>   sin_data_int <= to_unsigned(16339,N); cos_data_int <= to_unsigned(1205,N);
          when 977 =>   sin_data_int <= to_unsigned(16341,N); cos_data_int <= to_unsigned(1180,N);
          when 978 =>   sin_data_int <= to_unsigned(16343,N); cos_data_int <= to_unsigned(1155,N);
          when 979 =>   sin_data_int <= to_unsigned(16344,N); cos_data_int <= to_unsigned(1130,N);
          when 980 =>   sin_data_int <= to_unsigned(16346,N); cos_data_int <= to_unsigned(1105,N);
          when 981 =>   sin_data_int <= to_unsigned(16348,N); cos_data_int <= to_unsigned(1079,N);
          when 982 =>   sin_data_int <= to_unsigned(16350,N); cos_data_int <= to_unsigned(1054,N);
          when 983 =>   sin_data_int <= to_unsigned(16351,N); cos_data_int <= to_unsigned(1029,N);
          when 984 =>   sin_data_int <= to_unsigned(16353,N); cos_data_int <= to_unsigned(1004,N);
          when 985 =>   sin_data_int <= to_unsigned(16354,N); cos_data_int <= to_unsigned(979,N);
          when 986 =>   sin_data_int <= to_unsigned(16356,N); cos_data_int <= to_unsigned(954,N);
          when 987 =>   sin_data_int <= to_unsigned(16357,N); cos_data_int <= to_unsigned(929,N);
          when 988 =>   sin_data_int <= to_unsigned(16359,N); cos_data_int <= to_unsigned(904,N);
          when 989 =>   sin_data_int <= to_unsigned(16360,N); cos_data_int <= to_unsigned(879,N);
          when 990 =>   sin_data_int <= to_unsigned(16361,N); cos_data_int <= to_unsigned(854,N);
          when 991 =>   sin_data_int <= to_unsigned(16363,N); cos_data_int <= to_unsigned(829,N);
          when 992 =>   sin_data_int <= to_unsigned(16364,N); cos_data_int <= to_unsigned(803,N);
          when 993 =>   sin_data_int <= to_unsigned(16365,N); cos_data_int <= to_unsigned(778,N);
          when 994 =>   sin_data_int <= to_unsigned(16366,N); cos_data_int <= to_unsigned(753,N);
          when 995 =>   sin_data_int <= to_unsigned(16367,N); cos_data_int <= to_unsigned(728,N);
          when 996 =>   sin_data_int <= to_unsigned(16368,N); cos_data_int <= to_unsigned(703,N);
          when 997 =>   sin_data_int <= to_unsigned(16369,N); cos_data_int <= to_unsigned(678,N);
          when 998 =>   sin_data_int <= to_unsigned(16370,N); cos_data_int <= to_unsigned(653,N);
          when 999 =>   sin_data_int <= to_unsigned(16371,N); cos_data_int <= to_unsigned(628,N);
          when 1000 =>   sin_data_int <= to_unsigned(16372,N); cos_data_int <= to_unsigned(603,N);
          when 1001 =>   sin_data_int <= to_unsigned(16373,N); cos_data_int <= to_unsigned(577,N);
          when 1002 =>   sin_data_int <= to_unsigned(16374,N); cos_data_int <= to_unsigned(552,N);
          when 1003 =>   sin_data_int <= to_unsigned(16375,N); cos_data_int <= to_unsigned(527,N);
          when 1004 =>   sin_data_int <= to_unsigned(16376,N); cos_data_int <= to_unsigned(502,N);
          when 1005 =>   sin_data_int <= to_unsigned(16377,N); cos_data_int <= to_unsigned(477,N);
          when 1006 =>   sin_data_int <= to_unsigned(16377,N); cos_data_int <= to_unsigned(452,N);
          when 1007 =>   sin_data_int <= to_unsigned(16378,N); cos_data_int <= to_unsigned(427,N);
          when 1008 =>   sin_data_int <= to_unsigned(16379,N); cos_data_int <= to_unsigned(402,N);
          when 1009 =>   sin_data_int <= to_unsigned(16379,N); cos_data_int <= to_unsigned(376,N);
          when 1010 =>   sin_data_int <= to_unsigned(16380,N); cos_data_int <= to_unsigned(351,N);
          when 1011 =>   sin_data_int <= to_unsigned(16380,N); cos_data_int <= to_unsigned(326,N);
          when 1012 =>   sin_data_int <= to_unsigned(16381,N); cos_data_int <= to_unsigned(301,N);
          when 1013 =>   sin_data_int <= to_unsigned(16381,N); cos_data_int <= to_unsigned(276,N);
          when 1014 =>   sin_data_int <= to_unsigned(16382,N); cos_data_int <= to_unsigned(251,N);
          when 1015 =>   sin_data_int <= to_unsigned(16382,N); cos_data_int <= to_unsigned(226,N);
          when 1016 =>   sin_data_int <= to_unsigned(16382,N); cos_data_int <= to_unsigned(201,N);
          when 1017 =>   sin_data_int <= to_unsigned(16383,N); cos_data_int <= to_unsigned(175,N);
          when 1018 =>   sin_data_int <= to_unsigned(16383,N); cos_data_int <= to_unsigned(150,N);
          when 1019 =>   sin_data_int <= to_unsigned(16383,N); cos_data_int <= to_unsigned(125,N);
          when 1020 =>   sin_data_int <= to_unsigned(16383,N); cos_data_int <= to_unsigned(100,N);
          when 1021 =>   sin_data_int <= to_unsigned(16383,N); cos_data_int <= to_unsigned(75,N);
          when 1022 =>   sin_data_int <= to_unsigned(16383,N); cos_data_int <= to_unsigned(50,N);
          when 1023 =>   sin_data_int <= to_unsigned(16383,N); cos_data_int <= to_unsigned(25,N);
          when 1024 =>   sin_data_int <= to_unsigned(16384,N); cos_data_int <= to_unsigned(0,N);
          when 1025 =>   sin_data_int <= to_unsigned(16383,N); cos_data_int <= to_unsigned(65510,N);
          when 1026 =>   sin_data_int <= to_unsigned(16383,N); cos_data_int <= to_unsigned(65485,N);
          when 1027 =>   sin_data_int <= to_unsigned(16383,N); cos_data_int <= to_unsigned(65460,N);
          when 1028 =>   sin_data_int <= to_unsigned(16383,N); cos_data_int <= to_unsigned(65435,N);
          when 1029 =>   sin_data_int <= to_unsigned(16383,N); cos_data_int <= to_unsigned(65410,N);
          when 1030 =>   sin_data_int <= to_unsigned(16383,N); cos_data_int <= to_unsigned(65385,N);
          when 1031 =>   sin_data_int <= to_unsigned(16383,N); cos_data_int <= to_unsigned(65360,N);
          when 1032 =>   sin_data_int <= to_unsigned(16382,N); cos_data_int <= to_unsigned(65334,N);
          when 1033 =>   sin_data_int <= to_unsigned(16382,N); cos_data_int <= to_unsigned(65309,N);
          when 1034 =>   sin_data_int <= to_unsigned(16382,N); cos_data_int <= to_unsigned(65284,N);
          when 1035 =>   sin_data_int <= to_unsigned(16381,N); cos_data_int <= to_unsigned(65259,N);
          when 1036 =>   sin_data_int <= to_unsigned(16381,N); cos_data_int <= to_unsigned(65234,N);
          when 1037 =>   sin_data_int <= to_unsigned(16380,N); cos_data_int <= to_unsigned(65209,N);
          when 1038 =>   sin_data_int <= to_unsigned(16380,N); cos_data_int <= to_unsigned(65184,N);
          when 1039 =>   sin_data_int <= to_unsigned(16379,N); cos_data_int <= to_unsigned(65159,N);
          when 1040 =>   sin_data_int <= to_unsigned(16379,N); cos_data_int <= to_unsigned(65133,N);
          when 1041 =>   sin_data_int <= to_unsigned(16378,N); cos_data_int <= to_unsigned(65108,N);
          when 1042 =>   sin_data_int <= to_unsigned(16377,N); cos_data_int <= to_unsigned(65083,N);
          when 1043 =>   sin_data_int <= to_unsigned(16377,N); cos_data_int <= to_unsigned(65058,N);
          when 1044 =>   sin_data_int <= to_unsigned(16376,N); cos_data_int <= to_unsigned(65033,N);
          when 1045 =>   sin_data_int <= to_unsigned(16375,N); cos_data_int <= to_unsigned(65008,N);
          when 1046 =>   sin_data_int <= to_unsigned(16374,N); cos_data_int <= to_unsigned(64983,N);
          when 1047 =>   sin_data_int <= to_unsigned(16373,N); cos_data_int <= to_unsigned(64958,N);
          when 1048 =>   sin_data_int <= to_unsigned(16372,N); cos_data_int <= to_unsigned(64932,N);
          when 1049 =>   sin_data_int <= to_unsigned(16371,N); cos_data_int <= to_unsigned(64907,N);
          when 1050 =>   sin_data_int <= to_unsigned(16370,N); cos_data_int <= to_unsigned(64882,N);
          when 1051 =>   sin_data_int <= to_unsigned(16369,N); cos_data_int <= to_unsigned(64857,N);
          when 1052 =>   sin_data_int <= to_unsigned(16368,N); cos_data_int <= to_unsigned(64832,N);
          when 1053 =>   sin_data_int <= to_unsigned(16367,N); cos_data_int <= to_unsigned(64807,N);
          when 1054 =>   sin_data_int <= to_unsigned(16366,N); cos_data_int <= to_unsigned(64782,N);
          when 1055 =>   sin_data_int <= to_unsigned(16365,N); cos_data_int <= to_unsigned(64757,N);
          when 1056 =>   sin_data_int <= to_unsigned(16364,N); cos_data_int <= to_unsigned(64732,N);
          when 1057 =>   sin_data_int <= to_unsigned(16363,N); cos_data_int <= to_unsigned(64706,N);
          when 1058 =>   sin_data_int <= to_unsigned(16361,N); cos_data_int <= to_unsigned(64681,N);
          when 1059 =>   sin_data_int <= to_unsigned(16360,N); cos_data_int <= to_unsigned(64656,N);
          when 1060 =>   sin_data_int <= to_unsigned(16359,N); cos_data_int <= to_unsigned(64631,N);
          when 1061 =>   sin_data_int <= to_unsigned(16357,N); cos_data_int <= to_unsigned(64606,N);
          when 1062 =>   sin_data_int <= to_unsigned(16356,N); cos_data_int <= to_unsigned(64581,N);
          when 1063 =>   sin_data_int <= to_unsigned(16354,N); cos_data_int <= to_unsigned(64556,N);
          when 1064 =>   sin_data_int <= to_unsigned(16353,N); cos_data_int <= to_unsigned(64531,N);
          when 1065 =>   sin_data_int <= to_unsigned(16351,N); cos_data_int <= to_unsigned(64506,N);
          when 1066 =>   sin_data_int <= to_unsigned(16350,N); cos_data_int <= to_unsigned(64481,N);
          when 1067 =>   sin_data_int <= to_unsigned(16348,N); cos_data_int <= to_unsigned(64456,N);
          when 1068 =>   sin_data_int <= to_unsigned(16346,N); cos_data_int <= to_unsigned(64430,N);
          when 1069 =>   sin_data_int <= to_unsigned(16344,N); cos_data_int <= to_unsigned(64405,N);
          when 1070 =>   sin_data_int <= to_unsigned(16343,N); cos_data_int <= to_unsigned(64380,N);
          when 1071 =>   sin_data_int <= to_unsigned(16341,N); cos_data_int <= to_unsigned(64355,N);
          when 1072 =>   sin_data_int <= to_unsigned(16339,N); cos_data_int <= to_unsigned(64330,N);
          when 1073 =>   sin_data_int <= to_unsigned(16337,N); cos_data_int <= to_unsigned(64305,N);
          when 1074 =>   sin_data_int <= to_unsigned(16335,N); cos_data_int <= to_unsigned(64280,N);
          when 1075 =>   sin_data_int <= to_unsigned(16333,N); cos_data_int <= to_unsigned(64255,N);
          when 1076 =>   sin_data_int <= to_unsigned(16331,N); cos_data_int <= to_unsigned(64230,N);
          when 1077 =>   sin_data_int <= to_unsigned(16329,N); cos_data_int <= to_unsigned(64205,N);
          when 1078 =>   sin_data_int <= to_unsigned(16327,N); cos_data_int <= to_unsigned(64180,N);
          when 1079 =>   sin_data_int <= to_unsigned(16325,N); cos_data_int <= to_unsigned(64155,N);
          when 1080 =>   sin_data_int <= to_unsigned(16323,N); cos_data_int <= to_unsigned(64130,N);
          when 1081 =>   sin_data_int <= to_unsigned(16321,N); cos_data_int <= to_unsigned(64105,N);
          when 1082 =>   sin_data_int <= to_unsigned(16319,N); cos_data_int <= to_unsigned(64080,N);
          when 1083 =>   sin_data_int <= to_unsigned(16316,N); cos_data_int <= to_unsigned(64055,N);
          when 1084 =>   sin_data_int <= to_unsigned(16314,N); cos_data_int <= to_unsigned(64030,N);
          when 1085 =>   sin_data_int <= to_unsigned(16312,N); cos_data_int <= to_unsigned(64005,N);
          when 1086 =>   sin_data_int <= to_unsigned(16309,N); cos_data_int <= to_unsigned(63980,N);
          when 1087 =>   sin_data_int <= to_unsigned(16307,N); cos_data_int <= to_unsigned(63955,N);
          when 1088 =>   sin_data_int <= to_unsigned(16305,N); cos_data_int <= to_unsigned(63930,N);
          when 1089 =>   sin_data_int <= to_unsigned(16302,N); cos_data_int <= to_unsigned(63905,N);
          when 1090 =>   sin_data_int <= to_unsigned(16300,N); cos_data_int <= to_unsigned(63880,N);
          when 1091 =>   sin_data_int <= to_unsigned(16297,N); cos_data_int <= to_unsigned(63855,N);
          when 1092 =>   sin_data_int <= to_unsigned(16294,N); cos_data_int <= to_unsigned(63830,N);
          when 1093 =>   sin_data_int <= to_unsigned(16292,N); cos_data_int <= to_unsigned(63805,N);
          when 1094 =>   sin_data_int <= to_unsigned(16289,N); cos_data_int <= to_unsigned(63780,N);
          when 1095 =>   sin_data_int <= to_unsigned(16286,N); cos_data_int <= to_unsigned(63755,N);
          when 1096 =>   sin_data_int <= to_unsigned(16284,N); cos_data_int <= to_unsigned(63730,N);
          when 1097 =>   sin_data_int <= to_unsigned(16281,N); cos_data_int <= to_unsigned(63705,N);
          when 1098 =>   sin_data_int <= to_unsigned(16278,N); cos_data_int <= to_unsigned(63680,N);
          when 1099 =>   sin_data_int <= to_unsigned(16275,N); cos_data_int <= to_unsigned(63655,N);
          when 1100 =>   sin_data_int <= to_unsigned(16272,N); cos_data_int <= to_unsigned(63630,N);
          when 1101 =>   sin_data_int <= to_unsigned(16269,N); cos_data_int <= to_unsigned(63605,N);
          when 1102 =>   sin_data_int <= to_unsigned(16266,N); cos_data_int <= to_unsigned(63580,N);
          when 1103 =>   sin_data_int <= to_unsigned(16263,N); cos_data_int <= to_unsigned(63555,N);
          when 1104 =>   sin_data_int <= to_unsigned(16260,N); cos_data_int <= to_unsigned(63530,N);
          when 1105 =>   sin_data_int <= to_unsigned(16257,N); cos_data_int <= to_unsigned(63505,N);
          when 1106 =>   sin_data_int <= to_unsigned(16254,N); cos_data_int <= to_unsigned(63480,N);
          when 1107 =>   sin_data_int <= to_unsigned(16251,N); cos_data_int <= to_unsigned(63455,N);
          when 1108 =>   sin_data_int <= to_unsigned(16248,N); cos_data_int <= to_unsigned(63430,N);
          when 1109 =>   sin_data_int <= to_unsigned(16244,N); cos_data_int <= to_unsigned(63405,N);
          when 1110 =>   sin_data_int <= to_unsigned(16241,N); cos_data_int <= to_unsigned(63380,N);
          when 1111 =>   sin_data_int <= to_unsigned(16238,N); cos_data_int <= to_unsigned(63355,N);
          when 1112 =>   sin_data_int <= to_unsigned(16234,N); cos_data_int <= to_unsigned(63331,N);
          when 1113 =>   sin_data_int <= to_unsigned(16231,N); cos_data_int <= to_unsigned(63306,N);
          when 1114 =>   sin_data_int <= to_unsigned(16228,N); cos_data_int <= to_unsigned(63281,N);
          when 1115 =>   sin_data_int <= to_unsigned(16224,N); cos_data_int <= to_unsigned(63256,N);
          when 1116 =>   sin_data_int <= to_unsigned(16221,N); cos_data_int <= to_unsigned(63231,N);
          when 1117 =>   sin_data_int <= to_unsigned(16217,N); cos_data_int <= to_unsigned(63206,N);
          when 1118 =>   sin_data_int <= to_unsigned(16213,N); cos_data_int <= to_unsigned(63181,N);
          when 1119 =>   sin_data_int <= to_unsigned(16210,N); cos_data_int <= to_unsigned(63156,N);
          when 1120 =>   sin_data_int <= to_unsigned(16206,N); cos_data_int <= to_unsigned(63131,N);
          when 1121 =>   sin_data_int <= to_unsigned(16202,N); cos_data_int <= to_unsigned(63107,N);
          when 1122 =>   sin_data_int <= to_unsigned(16199,N); cos_data_int <= to_unsigned(63082,N);
          when 1123 =>   sin_data_int <= to_unsigned(16195,N); cos_data_int <= to_unsigned(63057,N);
          when 1124 =>   sin_data_int <= to_unsigned(16191,N); cos_data_int <= to_unsigned(63032,N);
          when 1125 =>   sin_data_int <= to_unsigned(16187,N); cos_data_int <= to_unsigned(63007,N);
          when 1126 =>   sin_data_int <= to_unsigned(16183,N); cos_data_int <= to_unsigned(62982,N);
          when 1127 =>   sin_data_int <= to_unsigned(16179,N); cos_data_int <= to_unsigned(62958,N);
          when 1128 =>   sin_data_int <= to_unsigned(16175,N); cos_data_int <= to_unsigned(62933,N);
          when 1129 =>   sin_data_int <= to_unsigned(16171,N); cos_data_int <= to_unsigned(62908,N);
          when 1130 =>   sin_data_int <= to_unsigned(16167,N); cos_data_int <= to_unsigned(62883,N);
          when 1131 =>   sin_data_int <= to_unsigned(16163,N); cos_data_int <= to_unsigned(62858,N);
          when 1132 =>   sin_data_int <= to_unsigned(16159,N); cos_data_int <= to_unsigned(62834,N);
          when 1133 =>   sin_data_int <= to_unsigned(16155,N); cos_data_int <= to_unsigned(62809,N);
          when 1134 =>   sin_data_int <= to_unsigned(16151,N); cos_data_int <= to_unsigned(62784,N);
          when 1135 =>   sin_data_int <= to_unsigned(16147,N); cos_data_int <= to_unsigned(62759,N);
          when 1136 =>   sin_data_int <= to_unsigned(16142,N); cos_data_int <= to_unsigned(62734,N);
          when 1137 =>   sin_data_int <= to_unsigned(16138,N); cos_data_int <= to_unsigned(62710,N);
          when 1138 =>   sin_data_int <= to_unsigned(16134,N); cos_data_int <= to_unsigned(62685,N);
          when 1139 =>   sin_data_int <= to_unsigned(16129,N); cos_data_int <= to_unsigned(62660,N);
          when 1140 =>   sin_data_int <= to_unsigned(16125,N); cos_data_int <= to_unsigned(62635,N);
          when 1141 =>   sin_data_int <= to_unsigned(16120,N); cos_data_int <= to_unsigned(62611,N);
          when 1142 =>   sin_data_int <= to_unsigned(16116,N); cos_data_int <= to_unsigned(62586,N);
          when 1143 =>   sin_data_int <= to_unsigned(16111,N); cos_data_int <= to_unsigned(62561,N);
          when 1144 =>   sin_data_int <= to_unsigned(16107,N); cos_data_int <= to_unsigned(62537,N);
          when 1145 =>   sin_data_int <= to_unsigned(16102,N); cos_data_int <= to_unsigned(62512,N);
          when 1146 =>   sin_data_int <= to_unsigned(16097,N); cos_data_int <= to_unsigned(62487,N);
          when 1147 =>   sin_data_int <= to_unsigned(16093,N); cos_data_int <= to_unsigned(62462,N);
          when 1148 =>   sin_data_int <= to_unsigned(16088,N); cos_data_int <= to_unsigned(62438,N);
          when 1149 =>   sin_data_int <= to_unsigned(16083,N); cos_data_int <= to_unsigned(62413,N);
          when 1150 =>   sin_data_int <= to_unsigned(16078,N); cos_data_int <= to_unsigned(62388,N);
          when 1151 =>   sin_data_int <= to_unsigned(16074,N); cos_data_int <= to_unsigned(62364,N);
          when 1152 =>   sin_data_int <= to_unsigned(16069,N); cos_data_int <= to_unsigned(62339,N);
          when 1153 =>   sin_data_int <= to_unsigned(16064,N); cos_data_int <= to_unsigned(62314,N);
          when 1154 =>   sin_data_int <= to_unsigned(16059,N); cos_data_int <= to_unsigned(62290,N);
          when 1155 =>   sin_data_int <= to_unsigned(16054,N); cos_data_int <= to_unsigned(62265,N);
          when 1156 =>   sin_data_int <= to_unsigned(16049,N); cos_data_int <= to_unsigned(62241,N);
          when 1157 =>   sin_data_int <= to_unsigned(16044,N); cos_data_int <= to_unsigned(62216,N);
          when 1158 =>   sin_data_int <= to_unsigned(16039,N); cos_data_int <= to_unsigned(62191,N);
          when 1159 =>   sin_data_int <= to_unsigned(16033,N); cos_data_int <= to_unsigned(62167,N);
          when 1160 =>   sin_data_int <= to_unsigned(16028,N); cos_data_int <= to_unsigned(62142,N);
          when 1161 =>   sin_data_int <= to_unsigned(16023,N); cos_data_int <= to_unsigned(62118,N);
          when 1162 =>   sin_data_int <= to_unsigned(16018,N); cos_data_int <= to_unsigned(62093,N);
          when 1163 =>   sin_data_int <= to_unsigned(16012,N); cos_data_int <= to_unsigned(62068,N);
          when 1164 =>   sin_data_int <= to_unsigned(16007,N); cos_data_int <= to_unsigned(62044,N);
          when 1165 =>   sin_data_int <= to_unsigned(16002,N); cos_data_int <= to_unsigned(62019,N);
          when 1166 =>   sin_data_int <= to_unsigned(15996,N); cos_data_int <= to_unsigned(61995,N);
          when 1167 =>   sin_data_int <= to_unsigned(15991,N); cos_data_int <= to_unsigned(61970,N);
          when 1168 =>   sin_data_int <= to_unsigned(15985,N); cos_data_int <= to_unsigned(61946,N);
          when 1169 =>   sin_data_int <= to_unsigned(15980,N); cos_data_int <= to_unsigned(61921,N);
          when 1170 =>   sin_data_int <= to_unsigned(15974,N); cos_data_int <= to_unsigned(61897,N);
          when 1171 =>   sin_data_int <= to_unsigned(15969,N); cos_data_int <= to_unsigned(61872,N);
          when 1172 =>   sin_data_int <= to_unsigned(15963,N); cos_data_int <= to_unsigned(61848,N);
          when 1173 =>   sin_data_int <= to_unsigned(15957,N); cos_data_int <= to_unsigned(61823,N);
          when 1174 =>   sin_data_int <= to_unsigned(15952,N); cos_data_int <= to_unsigned(61799,N);
          when 1175 =>   sin_data_int <= to_unsigned(15946,N); cos_data_int <= to_unsigned(61774,N);
          when 1176 =>   sin_data_int <= to_unsigned(15940,N); cos_data_int <= to_unsigned(61750,N);
          when 1177 =>   sin_data_int <= to_unsigned(15934,N); cos_data_int <= to_unsigned(61725,N);
          when 1178 =>   sin_data_int <= to_unsigned(15928,N); cos_data_int <= to_unsigned(61701,N);
          when 1179 =>   sin_data_int <= to_unsigned(15923,N); cos_data_int <= to_unsigned(61677,N);
          when 1180 =>   sin_data_int <= to_unsigned(15917,N); cos_data_int <= to_unsigned(61652,N);
          when 1181 =>   sin_data_int <= to_unsigned(15911,N); cos_data_int <= to_unsigned(61628,N);
          when 1182 =>   sin_data_int <= to_unsigned(15905,N); cos_data_int <= to_unsigned(61603,N);
          when 1183 =>   sin_data_int <= to_unsigned(15899,N); cos_data_int <= to_unsigned(61579,N);
          when 1184 =>   sin_data_int <= to_unsigned(15892,N); cos_data_int <= to_unsigned(61555,N);
          when 1185 =>   sin_data_int <= to_unsigned(15886,N); cos_data_int <= to_unsigned(61530,N);
          when 1186 =>   sin_data_int <= to_unsigned(15880,N); cos_data_int <= to_unsigned(61506,N);
          when 1187 =>   sin_data_int <= to_unsigned(15874,N); cos_data_int <= to_unsigned(61481,N);
          when 1188 =>   sin_data_int <= to_unsigned(15868,N); cos_data_int <= to_unsigned(61457,N);
          when 1189 =>   sin_data_int <= to_unsigned(15861,N); cos_data_int <= to_unsigned(61433,N);
          when 1190 =>   sin_data_int <= to_unsigned(15855,N); cos_data_int <= to_unsigned(61408,N);
          when 1191 =>   sin_data_int <= to_unsigned(15849,N); cos_data_int <= to_unsigned(61384,N);
          when 1192 =>   sin_data_int <= to_unsigned(15842,N); cos_data_int <= to_unsigned(61360,N);
          when 1193 =>   sin_data_int <= to_unsigned(15836,N); cos_data_int <= to_unsigned(61335,N);
          when 1194 =>   sin_data_int <= to_unsigned(15830,N); cos_data_int <= to_unsigned(61311,N);
          when 1195 =>   sin_data_int <= to_unsigned(15823,N); cos_data_int <= to_unsigned(61287,N);
          when 1196 =>   sin_data_int <= to_unsigned(15817,N); cos_data_int <= to_unsigned(61263,N);
          when 1197 =>   sin_data_int <= to_unsigned(15810,N); cos_data_int <= to_unsigned(61238,N);
          when 1198 =>   sin_data_int <= to_unsigned(15803,N); cos_data_int <= to_unsigned(61214,N);
          when 1199 =>   sin_data_int <= to_unsigned(15797,N); cos_data_int <= to_unsigned(61190,N);
          when 1200 =>   sin_data_int <= to_unsigned(15790,N); cos_data_int <= to_unsigned(61166,N);
          when 1201 =>   sin_data_int <= to_unsigned(15783,N); cos_data_int <= to_unsigned(61141,N);
          when 1202 =>   sin_data_int <= to_unsigned(15777,N); cos_data_int <= to_unsigned(61117,N);
          when 1203 =>   sin_data_int <= to_unsigned(15770,N); cos_data_int <= to_unsigned(61093,N);
          when 1204 =>   sin_data_int <= to_unsigned(15763,N); cos_data_int <= to_unsigned(61069,N);
          when 1205 =>   sin_data_int <= to_unsigned(15756,N); cos_data_int <= to_unsigned(61045,N);
          when 1206 =>   sin_data_int <= to_unsigned(15749,N); cos_data_int <= to_unsigned(61021,N);
          when 1207 =>   sin_data_int <= to_unsigned(15742,N); cos_data_int <= to_unsigned(60996,N);
          when 1208 =>   sin_data_int <= to_unsigned(15735,N); cos_data_int <= to_unsigned(60972,N);
          when 1209 =>   sin_data_int <= to_unsigned(15728,N); cos_data_int <= to_unsigned(60948,N);
          when 1210 =>   sin_data_int <= to_unsigned(15721,N); cos_data_int <= to_unsigned(60924,N);
          when 1211 =>   sin_data_int <= to_unsigned(15714,N); cos_data_int <= to_unsigned(60900,N);
          when 1212 =>   sin_data_int <= to_unsigned(15707,N); cos_data_int <= to_unsigned(60876,N);
          when 1213 =>   sin_data_int <= to_unsigned(15700,N); cos_data_int <= to_unsigned(60852,N);
          when 1214 =>   sin_data_int <= to_unsigned(15693,N); cos_data_int <= to_unsigned(60828,N);
          when 1215 =>   sin_data_int <= to_unsigned(15685,N); cos_data_int <= to_unsigned(60804,N);
          when 1216 =>   sin_data_int <= to_unsigned(15678,N); cos_data_int <= to_unsigned(60779,N);
          when 1217 =>   sin_data_int <= to_unsigned(15671,N); cos_data_int <= to_unsigned(60755,N);
          when 1218 =>   sin_data_int <= to_unsigned(15663,N); cos_data_int <= to_unsigned(60731,N);
          when 1219 =>   sin_data_int <= to_unsigned(15656,N); cos_data_int <= to_unsigned(60707,N);
          when 1220 =>   sin_data_int <= to_unsigned(15649,N); cos_data_int <= to_unsigned(60683,N);
          when 1221 =>   sin_data_int <= to_unsigned(15641,N); cos_data_int <= to_unsigned(60659,N);
          when 1222 =>   sin_data_int <= to_unsigned(15634,N); cos_data_int <= to_unsigned(60635,N);
          when 1223 =>   sin_data_int <= to_unsigned(15626,N); cos_data_int <= to_unsigned(60611,N);
          when 1224 =>   sin_data_int <= to_unsigned(15618,N); cos_data_int <= to_unsigned(60587,N);
          when 1225 =>   sin_data_int <= to_unsigned(15611,N); cos_data_int <= to_unsigned(60563,N);
          when 1226 =>   sin_data_int <= to_unsigned(15603,N); cos_data_int <= to_unsigned(60540,N);
          when 1227 =>   sin_data_int <= to_unsigned(15596,N); cos_data_int <= to_unsigned(60516,N);
          when 1228 =>   sin_data_int <= to_unsigned(15588,N); cos_data_int <= to_unsigned(60492,N);
          when 1229 =>   sin_data_int <= to_unsigned(15580,N); cos_data_int <= to_unsigned(60468,N);
          when 1230 =>   sin_data_int <= to_unsigned(15572,N); cos_data_int <= to_unsigned(60444,N);
          when 1231 =>   sin_data_int <= to_unsigned(15564,N); cos_data_int <= to_unsigned(60420,N);
          when 1232 =>   sin_data_int <= to_unsigned(15557,N); cos_data_int <= to_unsigned(60396,N);
          when 1233 =>   sin_data_int <= to_unsigned(15549,N); cos_data_int <= to_unsigned(60372,N);
          when 1234 =>   sin_data_int <= to_unsigned(15541,N); cos_data_int <= to_unsigned(60348,N);
          when 1235 =>   sin_data_int <= to_unsigned(15533,N); cos_data_int <= to_unsigned(60325,N);
          when 1236 =>   sin_data_int <= to_unsigned(15525,N); cos_data_int <= to_unsigned(60301,N);
          when 1237 =>   sin_data_int <= to_unsigned(15517,N); cos_data_int <= to_unsigned(60277,N);
          when 1238 =>   sin_data_int <= to_unsigned(15509,N); cos_data_int <= to_unsigned(60253,N);
          when 1239 =>   sin_data_int <= to_unsigned(15500,N); cos_data_int <= to_unsigned(60229,N);
          when 1240 =>   sin_data_int <= to_unsigned(15492,N); cos_data_int <= to_unsigned(60206,N);
          when 1241 =>   sin_data_int <= to_unsigned(15484,N); cos_data_int <= to_unsigned(60182,N);
          when 1242 =>   sin_data_int <= to_unsigned(15476,N); cos_data_int <= to_unsigned(60158,N);
          when 1243 =>   sin_data_int <= to_unsigned(15468,N); cos_data_int <= to_unsigned(60134,N);
          when 1244 =>   sin_data_int <= to_unsigned(15459,N); cos_data_int <= to_unsigned(60111,N);
          when 1245 =>   sin_data_int <= to_unsigned(15451,N); cos_data_int <= to_unsigned(60087,N);
          when 1246 =>   sin_data_int <= to_unsigned(15443,N); cos_data_int <= to_unsigned(60063,N);
          when 1247 =>   sin_data_int <= to_unsigned(15434,N); cos_data_int <= to_unsigned(60040,N);
          when 1248 =>   sin_data_int <= to_unsigned(15426,N); cos_data_int <= to_unsigned(60016,N);
          when 1249 =>   sin_data_int <= to_unsigned(15417,N); cos_data_int <= to_unsigned(59992,N);
          when 1250 =>   sin_data_int <= to_unsigned(15409,N); cos_data_int <= to_unsigned(59969,N);
          when 1251 =>   sin_data_int <= to_unsigned(15400,N); cos_data_int <= to_unsigned(59945,N);
          when 1252 =>   sin_data_int <= to_unsigned(15392,N); cos_data_int <= to_unsigned(59921,N);
          when 1253 =>   sin_data_int <= to_unsigned(15383,N); cos_data_int <= to_unsigned(59898,N);
          when 1254 =>   sin_data_int <= to_unsigned(15374,N); cos_data_int <= to_unsigned(59874,N);
          when 1255 =>   sin_data_int <= to_unsigned(15366,N); cos_data_int <= to_unsigned(59851,N);
          when 1256 =>   sin_data_int <= to_unsigned(15357,N); cos_data_int <= to_unsigned(59827,N);
          when 1257 =>   sin_data_int <= to_unsigned(15348,N); cos_data_int <= to_unsigned(59803,N);
          when 1258 =>   sin_data_int <= to_unsigned(15339,N); cos_data_int <= to_unsigned(59780,N);
          when 1259 =>   sin_data_int <= to_unsigned(15330,N); cos_data_int <= to_unsigned(59756,N);
          when 1260 =>   sin_data_int <= to_unsigned(15322,N); cos_data_int <= to_unsigned(59733,N);
          when 1261 =>   sin_data_int <= to_unsigned(15313,N); cos_data_int <= to_unsigned(59709,N);
          when 1262 =>   sin_data_int <= to_unsigned(15304,N); cos_data_int <= to_unsigned(59686,N);
          when 1263 =>   sin_data_int <= to_unsigned(15295,N); cos_data_int <= to_unsigned(59662,N);
          when 1264 =>   sin_data_int <= to_unsigned(15286,N); cos_data_int <= to_unsigned(59639,N);
          when 1265 =>   sin_data_int <= to_unsigned(15277,N); cos_data_int <= to_unsigned(59616,N);
          when 1266 =>   sin_data_int <= to_unsigned(15267,N); cos_data_int <= to_unsigned(59592,N);
          when 1267 =>   sin_data_int <= to_unsigned(15258,N); cos_data_int <= to_unsigned(59569,N);
          when 1268 =>   sin_data_int <= to_unsigned(15249,N); cos_data_int <= to_unsigned(59545,N);
          when 1269 =>   sin_data_int <= to_unsigned(15240,N); cos_data_int <= to_unsigned(59522,N);
          when 1270 =>   sin_data_int <= to_unsigned(15231,N); cos_data_int <= to_unsigned(59499,N);
          when 1271 =>   sin_data_int <= to_unsigned(15221,N); cos_data_int <= to_unsigned(59475,N);
          when 1272 =>   sin_data_int <= to_unsigned(15212,N); cos_data_int <= to_unsigned(59452,N);
          when 1273 =>   sin_data_int <= to_unsigned(15203,N); cos_data_int <= to_unsigned(59429,N);
          when 1274 =>   sin_data_int <= to_unsigned(15193,N); cos_data_int <= to_unsigned(59405,N);
          when 1275 =>   sin_data_int <= to_unsigned(15184,N); cos_data_int <= to_unsigned(59382,N);
          when 1276 =>   sin_data_int <= to_unsigned(15175,N); cos_data_int <= to_unsigned(59359,N);
          when 1277 =>   sin_data_int <= to_unsigned(15165,N); cos_data_int <= to_unsigned(59335,N);
          when 1278 =>   sin_data_int <= to_unsigned(15156,N); cos_data_int <= to_unsigned(59312,N);
          when 1279 =>   sin_data_int <= to_unsigned(15146,N); cos_data_int <= to_unsigned(59289,N);
          when 1280 =>   sin_data_int <= to_unsigned(15136,N); cos_data_int <= to_unsigned(59266,N);
          when 1281 =>   sin_data_int <= to_unsigned(15127,N); cos_data_int <= to_unsigned(59242,N);
          when 1282 =>   sin_data_int <= to_unsigned(15117,N); cos_data_int <= to_unsigned(59219,N);
          when 1283 =>   sin_data_int <= to_unsigned(15107,N); cos_data_int <= to_unsigned(59196,N);
          when 1284 =>   sin_data_int <= to_unsigned(15098,N); cos_data_int <= to_unsigned(59173,N);
          when 1285 =>   sin_data_int <= to_unsigned(15088,N); cos_data_int <= to_unsigned(59150,N);
          when 1286 =>   sin_data_int <= to_unsigned(15078,N); cos_data_int <= to_unsigned(59127,N);
          when 1287 =>   sin_data_int <= to_unsigned(15068,N); cos_data_int <= to_unsigned(59103,N);
          when 1288 =>   sin_data_int <= to_unsigned(15058,N); cos_data_int <= to_unsigned(59080,N);
          when 1289 =>   sin_data_int <= to_unsigned(15048,N); cos_data_int <= to_unsigned(59057,N);
          when 1290 =>   sin_data_int <= to_unsigned(15038,N); cos_data_int <= to_unsigned(59034,N);
          when 1291 =>   sin_data_int <= to_unsigned(15028,N); cos_data_int <= to_unsigned(59011,N);
          when 1292 =>   sin_data_int <= to_unsigned(15018,N); cos_data_int <= to_unsigned(58988,N);
          when 1293 =>   sin_data_int <= to_unsigned(15008,N); cos_data_int <= to_unsigned(58965,N);
          when 1294 =>   sin_data_int <= to_unsigned(14998,N); cos_data_int <= to_unsigned(58942,N);
          when 1295 =>   sin_data_int <= to_unsigned(14988,N); cos_data_int <= to_unsigned(58919,N);
          when 1296 =>   sin_data_int <= to_unsigned(14978,N); cos_data_int <= to_unsigned(58896,N);
          when 1297 =>   sin_data_int <= to_unsigned(14968,N); cos_data_int <= to_unsigned(58873,N);
          when 1298 =>   sin_data_int <= to_unsigned(14957,N); cos_data_int <= to_unsigned(58850,N);
          when 1299 =>   sin_data_int <= to_unsigned(14947,N); cos_data_int <= to_unsigned(58827,N);
          when 1300 =>   sin_data_int <= to_unsigned(14937,N); cos_data_int <= to_unsigned(58804,N);
          when 1301 =>   sin_data_int <= to_unsigned(14927,N); cos_data_int <= to_unsigned(58781,N);
          when 1302 =>   sin_data_int <= to_unsigned(14916,N); cos_data_int <= to_unsigned(58758,N);
          when 1303 =>   sin_data_int <= to_unsigned(14906,N); cos_data_int <= to_unsigned(58736,N);
          when 1304 =>   sin_data_int <= to_unsigned(14895,N); cos_data_int <= to_unsigned(58713,N);
          when 1305 =>   sin_data_int <= to_unsigned(14885,N); cos_data_int <= to_unsigned(58690,N);
          when 1306 =>   sin_data_int <= to_unsigned(14874,N); cos_data_int <= to_unsigned(58667,N);
          when 1307 =>   sin_data_int <= to_unsigned(14864,N); cos_data_int <= to_unsigned(58644,N);
          when 1308 =>   sin_data_int <= to_unsigned(14853,N); cos_data_int <= to_unsigned(58621,N);
          when 1309 =>   sin_data_int <= to_unsigned(14843,N); cos_data_int <= to_unsigned(58599,N);
          when 1310 =>   sin_data_int <= to_unsigned(14832,N); cos_data_int <= to_unsigned(58576,N);
          when 1311 =>   sin_data_int <= to_unsigned(14821,N); cos_data_int <= to_unsigned(58553,N);
          when 1312 =>   sin_data_int <= to_unsigned(14810,N); cos_data_int <= to_unsigned(58530,N);
          when 1313 =>   sin_data_int <= to_unsigned(14800,N); cos_data_int <= to_unsigned(58508,N);
          when 1314 =>   sin_data_int <= to_unsigned(14789,N); cos_data_int <= to_unsigned(58485,N);
          when 1315 =>   sin_data_int <= to_unsigned(14778,N); cos_data_int <= to_unsigned(58462,N);
          when 1316 =>   sin_data_int <= to_unsigned(14767,N); cos_data_int <= to_unsigned(58440,N);
          when 1317 =>   sin_data_int <= to_unsigned(14756,N); cos_data_int <= to_unsigned(58417,N);
          when 1318 =>   sin_data_int <= to_unsigned(14745,N); cos_data_int <= to_unsigned(58394,N);
          when 1319 =>   sin_data_int <= to_unsigned(14734,N); cos_data_int <= to_unsigned(58372,N);
          when 1320 =>   sin_data_int <= to_unsigned(14723,N); cos_data_int <= to_unsigned(58349,N);
          when 1321 =>   sin_data_int <= to_unsigned(14712,N); cos_data_int <= to_unsigned(58327,N);
          when 1322 =>   sin_data_int <= to_unsigned(14701,N); cos_data_int <= to_unsigned(58304,N);
          when 1323 =>   sin_data_int <= to_unsigned(14690,N); cos_data_int <= to_unsigned(58282,N);
          when 1324 =>   sin_data_int <= to_unsigned(14679,N); cos_data_int <= to_unsigned(58259,N);
          when 1325 =>   sin_data_int <= to_unsigned(14668,N); cos_data_int <= to_unsigned(58236,N);
          when 1326 =>   sin_data_int <= to_unsigned(14657,N); cos_data_int <= to_unsigned(58214,N);
          when 1327 =>   sin_data_int <= to_unsigned(14645,N); cos_data_int <= to_unsigned(58192,N);
          when 1328 =>   sin_data_int <= to_unsigned(14634,N); cos_data_int <= to_unsigned(58169,N);
          when 1329 =>   sin_data_int <= to_unsigned(14623,N); cos_data_int <= to_unsigned(58147,N);
          when 1330 =>   sin_data_int <= to_unsigned(14611,N); cos_data_int <= to_unsigned(58124,N);
          when 1331 =>   sin_data_int <= to_unsigned(14600,N); cos_data_int <= to_unsigned(58102,N);
          when 1332 =>   sin_data_int <= to_unsigned(14589,N); cos_data_int <= to_unsigned(58079,N);
          when 1333 =>   sin_data_int <= to_unsigned(14577,N); cos_data_int <= to_unsigned(58057,N);
          when 1334 =>   sin_data_int <= to_unsigned(14566,N); cos_data_int <= to_unsigned(58035,N);
          when 1335 =>   sin_data_int <= to_unsigned(14554,N); cos_data_int <= to_unsigned(58012,N);
          when 1336 =>   sin_data_int <= to_unsigned(14543,N); cos_data_int <= to_unsigned(57990,N);
          when 1337 =>   sin_data_int <= to_unsigned(14531,N); cos_data_int <= to_unsigned(57968,N);
          when 1338 =>   sin_data_int <= to_unsigned(14519,N); cos_data_int <= to_unsigned(57945,N);
          when 1339 =>   sin_data_int <= to_unsigned(14508,N); cos_data_int <= to_unsigned(57923,N);
          when 1340 =>   sin_data_int <= to_unsigned(14496,N); cos_data_int <= to_unsigned(57901,N);
          when 1341 =>   sin_data_int <= to_unsigned(14484,N); cos_data_int <= to_unsigned(57879,N);
          when 1342 =>   sin_data_int <= to_unsigned(14473,N); cos_data_int <= to_unsigned(57857,N);
          when 1343 =>   sin_data_int <= to_unsigned(14461,N); cos_data_int <= to_unsigned(57834,N);
          when 1344 =>   sin_data_int <= to_unsigned(14449,N); cos_data_int <= to_unsigned(57812,N);
          when 1345 =>   sin_data_int <= to_unsigned(14437,N); cos_data_int <= to_unsigned(57790,N);
          when 1346 =>   sin_data_int <= to_unsigned(14425,N); cos_data_int <= to_unsigned(57768,N);
          when 1347 =>   sin_data_int <= to_unsigned(14413,N); cos_data_int <= to_unsigned(57746,N);
          when 1348 =>   sin_data_int <= to_unsigned(14401,N); cos_data_int <= to_unsigned(57724,N);
          when 1349 =>   sin_data_int <= to_unsigned(14389,N); cos_data_int <= to_unsigned(57702,N);
          when 1350 =>   sin_data_int <= to_unsigned(14377,N); cos_data_int <= to_unsigned(57679,N);
          when 1351 =>   sin_data_int <= to_unsigned(14365,N); cos_data_int <= to_unsigned(57657,N);
          when 1352 =>   sin_data_int <= to_unsigned(14353,N); cos_data_int <= to_unsigned(57635,N);
          when 1353 =>   sin_data_int <= to_unsigned(14341,N); cos_data_int <= to_unsigned(57613,N);
          when 1354 =>   sin_data_int <= to_unsigned(14329,N); cos_data_int <= to_unsigned(57591,N);
          when 1355 =>   sin_data_int <= to_unsigned(14317,N); cos_data_int <= to_unsigned(57569,N);
          when 1356 =>   sin_data_int <= to_unsigned(14304,N); cos_data_int <= to_unsigned(57547,N);
          when 1357 =>   sin_data_int <= to_unsigned(14292,N); cos_data_int <= to_unsigned(57526,N);
          when 1358 =>   sin_data_int <= to_unsigned(14280,N); cos_data_int <= to_unsigned(57504,N);
          when 1359 =>   sin_data_int <= to_unsigned(14267,N); cos_data_int <= to_unsigned(57482,N);
          when 1360 =>   sin_data_int <= to_unsigned(14255,N); cos_data_int <= to_unsigned(57460,N);
          when 1361 =>   sin_data_int <= to_unsigned(14243,N); cos_data_int <= to_unsigned(57438,N);
          when 1362 =>   sin_data_int <= to_unsigned(14230,N); cos_data_int <= to_unsigned(57416,N);
          when 1363 =>   sin_data_int <= to_unsigned(14218,N); cos_data_int <= to_unsigned(57394,N);
          when 1364 =>   sin_data_int <= to_unsigned(14205,N); cos_data_int <= to_unsigned(57373,N);
          when 1365 =>   sin_data_int <= to_unsigned(14193,N); cos_data_int <= to_unsigned(57351,N);
          when 1366 =>   sin_data_int <= to_unsigned(14180,N); cos_data_int <= to_unsigned(57329,N);
          when 1367 =>   sin_data_int <= to_unsigned(14167,N); cos_data_int <= to_unsigned(57307,N);
          when 1368 =>   sin_data_int <= to_unsigned(14155,N); cos_data_int <= to_unsigned(57286,N);
          when 1369 =>   sin_data_int <= to_unsigned(14142,N); cos_data_int <= to_unsigned(57264,N);
          when 1370 =>   sin_data_int <= to_unsigned(14129,N); cos_data_int <= to_unsigned(57242,N);
          when 1371 =>   sin_data_int <= to_unsigned(14117,N); cos_data_int <= to_unsigned(57220,N);
          when 1372 =>   sin_data_int <= to_unsigned(14104,N); cos_data_int <= to_unsigned(57199,N);
          when 1373 =>   sin_data_int <= to_unsigned(14091,N); cos_data_int <= to_unsigned(57177,N);
          when 1374 =>   sin_data_int <= to_unsigned(14078,N); cos_data_int <= to_unsigned(57156,N);
          when 1375 =>   sin_data_int <= to_unsigned(14065,N); cos_data_int <= to_unsigned(57134,N);
          when 1376 =>   sin_data_int <= to_unsigned(14053,N); cos_data_int <= to_unsigned(57112,N);
          when 1377 =>   sin_data_int <= to_unsigned(14040,N); cos_data_int <= to_unsigned(57091,N);
          when 1378 =>   sin_data_int <= to_unsigned(14027,N); cos_data_int <= to_unsigned(57069,N);
          when 1379 =>   sin_data_int <= to_unsigned(14014,N); cos_data_int <= to_unsigned(57048,N);
          when 1380 =>   sin_data_int <= to_unsigned(14001,N); cos_data_int <= to_unsigned(57026,N);
          when 1381 =>   sin_data_int <= to_unsigned(13988,N); cos_data_int <= to_unsigned(57005,N);
          when 1382 =>   sin_data_int <= to_unsigned(13974,N); cos_data_int <= to_unsigned(56983,N);
          when 1383 =>   sin_data_int <= to_unsigned(13961,N); cos_data_int <= to_unsigned(56962,N);
          when 1384 =>   sin_data_int <= to_unsigned(13948,N); cos_data_int <= to_unsigned(56941,N);
          when 1385 =>   sin_data_int <= to_unsigned(13935,N); cos_data_int <= to_unsigned(56919,N);
          when 1386 =>   sin_data_int <= to_unsigned(13922,N); cos_data_int <= to_unsigned(56898,N);
          when 1387 =>   sin_data_int <= to_unsigned(13908,N); cos_data_int <= to_unsigned(56877,N);
          when 1388 =>   sin_data_int <= to_unsigned(13895,N); cos_data_int <= to_unsigned(56855,N);
          when 1389 =>   sin_data_int <= to_unsigned(13882,N); cos_data_int <= to_unsigned(56834,N);
          when 1390 =>   sin_data_int <= to_unsigned(13868,N); cos_data_int <= to_unsigned(56813,N);
          when 1391 =>   sin_data_int <= to_unsigned(13855,N); cos_data_int <= to_unsigned(56791,N);
          when 1392 =>   sin_data_int <= to_unsigned(13842,N); cos_data_int <= to_unsigned(56770,N);
          when 1393 =>   sin_data_int <= to_unsigned(13828,N); cos_data_int <= to_unsigned(56749,N);
          when 1394 =>   sin_data_int <= to_unsigned(13815,N); cos_data_int <= to_unsigned(56728,N);
          when 1395 =>   sin_data_int <= to_unsigned(13801,N); cos_data_int <= to_unsigned(56706,N);
          when 1396 =>   sin_data_int <= to_unsigned(13788,N); cos_data_int <= to_unsigned(56685,N);
          when 1397 =>   sin_data_int <= to_unsigned(13774,N); cos_data_int <= to_unsigned(56664,N);
          when 1398 =>   sin_data_int <= to_unsigned(13760,N); cos_data_int <= to_unsigned(56643,N);
          when 1399 =>   sin_data_int <= to_unsigned(13747,N); cos_data_int <= to_unsigned(56622,N);
          when 1400 =>   sin_data_int <= to_unsigned(13733,N); cos_data_int <= to_unsigned(56601,N);
          when 1401 =>   sin_data_int <= to_unsigned(13719,N); cos_data_int <= to_unsigned(56580,N);
          when 1402 =>   sin_data_int <= to_unsigned(13705,N); cos_data_int <= to_unsigned(56559,N);
          when 1403 =>   sin_data_int <= to_unsigned(13692,N); cos_data_int <= to_unsigned(56538,N);
          when 1404 =>   sin_data_int <= to_unsigned(13678,N); cos_data_int <= to_unsigned(56517,N);
          when 1405 =>   sin_data_int <= to_unsigned(13664,N); cos_data_int <= to_unsigned(56496,N);
          when 1406 =>   sin_data_int <= to_unsigned(13650,N); cos_data_int <= to_unsigned(56475,N);
          when 1407 =>   sin_data_int <= to_unsigned(13636,N); cos_data_int <= to_unsigned(56454,N);
          when 1408 =>   sin_data_int <= to_unsigned(13622,N); cos_data_int <= to_unsigned(56433,N);
          when 1409 =>   sin_data_int <= to_unsigned(13608,N); cos_data_int <= to_unsigned(56412,N);
          when 1410 =>   sin_data_int <= to_unsigned(13594,N); cos_data_int <= to_unsigned(56391,N);
          when 1411 =>   sin_data_int <= to_unsigned(13580,N); cos_data_int <= to_unsigned(56370,N);
          when 1412 =>   sin_data_int <= to_unsigned(13566,N); cos_data_int <= to_unsigned(56350,N);
          when 1413 =>   sin_data_int <= to_unsigned(13552,N); cos_data_int <= to_unsigned(56329,N);
          when 1414 =>   sin_data_int <= to_unsigned(13538,N); cos_data_int <= to_unsigned(56308,N);
          when 1415 =>   sin_data_int <= to_unsigned(13524,N); cos_data_int <= to_unsigned(56287,N);
          when 1416 =>   sin_data_int <= to_unsigned(13510,N); cos_data_int <= to_unsigned(56267,N);
          when 1417 =>   sin_data_int <= to_unsigned(13495,N); cos_data_int <= to_unsigned(56246,N);
          when 1418 =>   sin_data_int <= to_unsigned(13481,N); cos_data_int <= to_unsigned(56225,N);
          when 1419 =>   sin_data_int <= to_unsigned(13467,N); cos_data_int <= to_unsigned(56204,N);
          when 1420 =>   sin_data_int <= to_unsigned(13452,N); cos_data_int <= to_unsigned(56184,N);
          when 1421 =>   sin_data_int <= to_unsigned(13438,N); cos_data_int <= to_unsigned(56163,N);
          when 1422 =>   sin_data_int <= to_unsigned(13424,N); cos_data_int <= to_unsigned(56143,N);
          when 1423 =>   sin_data_int <= to_unsigned(13409,N); cos_data_int <= to_unsigned(56122,N);
          when 1424 =>   sin_data_int <= to_unsigned(13395,N); cos_data_int <= to_unsigned(56101,N);
          when 1425 =>   sin_data_int <= to_unsigned(13380,N); cos_data_int <= to_unsigned(56081,N);
          when 1426 =>   sin_data_int <= to_unsigned(13366,N); cos_data_int <= to_unsigned(56060,N);
          when 1427 =>   sin_data_int <= to_unsigned(13351,N); cos_data_int <= to_unsigned(56040,N);
          when 1428 =>   sin_data_int <= to_unsigned(13337,N); cos_data_int <= to_unsigned(56019,N);
          when 1429 =>   sin_data_int <= to_unsigned(13322,N); cos_data_int <= to_unsigned(55999,N);
          when 1430 =>   sin_data_int <= to_unsigned(13307,N); cos_data_int <= to_unsigned(55979,N);
          when 1431 =>   sin_data_int <= to_unsigned(13293,N); cos_data_int <= to_unsigned(55958,N);
          when 1432 =>   sin_data_int <= to_unsigned(13278,N); cos_data_int <= to_unsigned(55938,N);
          when 1433 =>   sin_data_int <= to_unsigned(13263,N); cos_data_int <= to_unsigned(55917,N);
          when 1434 =>   sin_data_int <= to_unsigned(13249,N); cos_data_int <= to_unsigned(55897,N);
          when 1435 =>   sin_data_int <= to_unsigned(13234,N); cos_data_int <= to_unsigned(55877,N);
          when 1436 =>   sin_data_int <= to_unsigned(13219,N); cos_data_int <= to_unsigned(55856,N);
          when 1437 =>   sin_data_int <= to_unsigned(13204,N); cos_data_int <= to_unsigned(55836,N);
          when 1438 =>   sin_data_int <= to_unsigned(13189,N); cos_data_int <= to_unsigned(55816,N);
          when 1439 =>   sin_data_int <= to_unsigned(13174,N); cos_data_int <= to_unsigned(55796,N);
          when 1440 =>   sin_data_int <= to_unsigned(13159,N); cos_data_int <= to_unsigned(55776,N);
          when 1441 =>   sin_data_int <= to_unsigned(13144,N); cos_data_int <= to_unsigned(55755,N);
          when 1442 =>   sin_data_int <= to_unsigned(13129,N); cos_data_int <= to_unsigned(55735,N);
          when 1443 =>   sin_data_int <= to_unsigned(13114,N); cos_data_int <= to_unsigned(55715,N);
          when 1444 =>   sin_data_int <= to_unsigned(13099,N); cos_data_int <= to_unsigned(55695,N);
          when 1445 =>   sin_data_int <= to_unsigned(13084,N); cos_data_int <= to_unsigned(55675,N);
          when 1446 =>   sin_data_int <= to_unsigned(13069,N); cos_data_int <= to_unsigned(55655,N);
          when 1447 =>   sin_data_int <= to_unsigned(13054,N); cos_data_int <= to_unsigned(55635,N);
          when 1448 =>   sin_data_int <= to_unsigned(13038,N); cos_data_int <= to_unsigned(55615,N);
          when 1449 =>   sin_data_int <= to_unsigned(13023,N); cos_data_int <= to_unsigned(55595,N);
          when 1450 =>   sin_data_int <= to_unsigned(13008,N); cos_data_int <= to_unsigned(55575,N);
          when 1451 =>   sin_data_int <= to_unsigned(12993,N); cos_data_int <= to_unsigned(55555,N);
          when 1452 =>   sin_data_int <= to_unsigned(12977,N); cos_data_int <= to_unsigned(55535,N);
          when 1453 =>   sin_data_int <= to_unsigned(12962,N); cos_data_int <= to_unsigned(55515,N);
          when 1454 =>   sin_data_int <= to_unsigned(12947,N); cos_data_int <= to_unsigned(55495,N);
          when 1455 =>   sin_data_int <= to_unsigned(12931,N); cos_data_int <= to_unsigned(55475,N);
          when 1456 =>   sin_data_int <= to_unsigned(12916,N); cos_data_int <= to_unsigned(55456,N);
          when 1457 =>   sin_data_int <= to_unsigned(12900,N); cos_data_int <= to_unsigned(55436,N);
          when 1458 =>   sin_data_int <= to_unsigned(12885,N); cos_data_int <= to_unsigned(55416,N);
          when 1459 =>   sin_data_int <= to_unsigned(12869,N); cos_data_int <= to_unsigned(55396,N);
          when 1460 =>   sin_data_int <= to_unsigned(12854,N); cos_data_int <= to_unsigned(55376,N);
          when 1461 =>   sin_data_int <= to_unsigned(12838,N); cos_data_int <= to_unsigned(55357,N);
          when 1462 =>   sin_data_int <= to_unsigned(12822,N); cos_data_int <= to_unsigned(55337,N);
          when 1463 =>   sin_data_int <= to_unsigned(12807,N); cos_data_int <= to_unsigned(55317,N);
          when 1464 =>   sin_data_int <= to_unsigned(12791,N); cos_data_int <= to_unsigned(55298,N);
          when 1465 =>   sin_data_int <= to_unsigned(12775,N); cos_data_int <= to_unsigned(55278,N);
          when 1466 =>   sin_data_int <= to_unsigned(12760,N); cos_data_int <= to_unsigned(55259,N);
          when 1467 =>   sin_data_int <= to_unsigned(12744,N); cos_data_int <= to_unsigned(55239,N);
          when 1468 =>   sin_data_int <= to_unsigned(12728,N); cos_data_int <= to_unsigned(55220,N);
          when 1469 =>   sin_data_int <= to_unsigned(12712,N); cos_data_int <= to_unsigned(55200,N);
          when 1470 =>   sin_data_int <= to_unsigned(12696,N); cos_data_int <= to_unsigned(55181,N);
          when 1471 =>   sin_data_int <= to_unsigned(12680,N); cos_data_int <= to_unsigned(55161,N);
          when 1472 =>   sin_data_int <= to_unsigned(12665,N); cos_data_int <= to_unsigned(55142,N);
          when 1473 =>   sin_data_int <= to_unsigned(12649,N); cos_data_int <= to_unsigned(55122,N);
          when 1474 =>   sin_data_int <= to_unsigned(12633,N); cos_data_int <= to_unsigned(55103,N);
          when 1475 =>   sin_data_int <= to_unsigned(12617,N); cos_data_int <= to_unsigned(55083,N);
          when 1476 =>   sin_data_int <= to_unsigned(12600,N); cos_data_int <= to_unsigned(55064,N);
          when 1477 =>   sin_data_int <= to_unsigned(12584,N); cos_data_int <= to_unsigned(55045,N);
          when 1478 =>   sin_data_int <= to_unsigned(12568,N); cos_data_int <= to_unsigned(55025,N);
          when 1479 =>   sin_data_int <= to_unsigned(12552,N); cos_data_int <= to_unsigned(55006,N);
          when 1480 =>   sin_data_int <= to_unsigned(12536,N); cos_data_int <= to_unsigned(54987,N);
          when 1481 =>   sin_data_int <= to_unsigned(12520,N); cos_data_int <= to_unsigned(54968,N);
          when 1482 =>   sin_data_int <= to_unsigned(12504,N); cos_data_int <= to_unsigned(54949,N);
          when 1483 =>   sin_data_int <= to_unsigned(12487,N); cos_data_int <= to_unsigned(54929,N);
          when 1484 =>   sin_data_int <= to_unsigned(12471,N); cos_data_int <= to_unsigned(54910,N);
          when 1485 =>   sin_data_int <= to_unsigned(12455,N); cos_data_int <= to_unsigned(54891,N);
          when 1486 =>   sin_data_int <= to_unsigned(12438,N); cos_data_int <= to_unsigned(54872,N);
          when 1487 =>   sin_data_int <= to_unsigned(12422,N); cos_data_int <= to_unsigned(54853,N);
          when 1488 =>   sin_data_int <= to_unsigned(12406,N); cos_data_int <= to_unsigned(54834,N);
          when 1489 =>   sin_data_int <= to_unsigned(12389,N); cos_data_int <= to_unsigned(54815,N);
          when 1490 =>   sin_data_int <= to_unsigned(12373,N); cos_data_int <= to_unsigned(54796,N);
          when 1491 =>   sin_data_int <= to_unsigned(12356,N); cos_data_int <= to_unsigned(54777,N);
          when 1492 =>   sin_data_int <= to_unsigned(12340,N); cos_data_int <= to_unsigned(54758,N);
          when 1493 =>   sin_data_int <= to_unsigned(12323,N); cos_data_int <= to_unsigned(54739,N);
          when 1494 =>   sin_data_int <= to_unsigned(12307,N); cos_data_int <= to_unsigned(54720,N);
          when 1495 =>   sin_data_int <= to_unsigned(12290,N); cos_data_int <= to_unsigned(54701,N);
          when 1496 =>   sin_data_int <= to_unsigned(12273,N); cos_data_int <= to_unsigned(54682,N);
          when 1497 =>   sin_data_int <= to_unsigned(12257,N); cos_data_int <= to_unsigned(54664,N);
          when 1498 =>   sin_data_int <= to_unsigned(12240,N); cos_data_int <= to_unsigned(54645,N);
          when 1499 =>   sin_data_int <= to_unsigned(12223,N); cos_data_int <= to_unsigned(54626,N);
          when 1500 =>   sin_data_int <= to_unsigned(12207,N); cos_data_int <= to_unsigned(54607,N);
          when 1501 =>   sin_data_int <= to_unsigned(12190,N); cos_data_int <= to_unsigned(54589,N);
          when 1502 =>   sin_data_int <= to_unsigned(12173,N); cos_data_int <= to_unsigned(54570,N);
          when 1503 =>   sin_data_int <= to_unsigned(12156,N); cos_data_int <= to_unsigned(54551,N);
          when 1504 =>   sin_data_int <= to_unsigned(12139,N); cos_data_int <= to_unsigned(54533,N);
          when 1505 =>   sin_data_int <= to_unsigned(12122,N); cos_data_int <= to_unsigned(54514,N);
          when 1506 =>   sin_data_int <= to_unsigned(12105,N); cos_data_int <= to_unsigned(54495,N);
          when 1507 =>   sin_data_int <= to_unsigned(12088,N); cos_data_int <= to_unsigned(54477,N);
          when 1508 =>   sin_data_int <= to_unsigned(12072,N); cos_data_int <= to_unsigned(54458,N);
          when 1509 =>   sin_data_int <= to_unsigned(12054,N); cos_data_int <= to_unsigned(54440,N);
          when 1510 =>   sin_data_int <= to_unsigned(12037,N); cos_data_int <= to_unsigned(54421,N);
          when 1511 =>   sin_data_int <= to_unsigned(12020,N); cos_data_int <= to_unsigned(54403,N);
          when 1512 =>   sin_data_int <= to_unsigned(12003,N); cos_data_int <= to_unsigned(54385,N);
          when 1513 =>   sin_data_int <= to_unsigned(11986,N); cos_data_int <= to_unsigned(54366,N);
          when 1514 =>   sin_data_int <= to_unsigned(11969,N); cos_data_int <= to_unsigned(54348,N);
          when 1515 =>   sin_data_int <= to_unsigned(11952,N); cos_data_int <= to_unsigned(54329,N);
          when 1516 =>   sin_data_int <= to_unsigned(11935,N); cos_data_int <= to_unsigned(54311,N);
          when 1517 =>   sin_data_int <= to_unsigned(11917,N); cos_data_int <= to_unsigned(54293,N);
          when 1518 =>   sin_data_int <= to_unsigned(11900,N); cos_data_int <= to_unsigned(54275,N);
          when 1519 =>   sin_data_int <= to_unsigned(11883,N); cos_data_int <= to_unsigned(54256,N);
          when 1520 =>   sin_data_int <= to_unsigned(11866,N); cos_data_int <= to_unsigned(54238,N);
          when 1521 =>   sin_data_int <= to_unsigned(11848,N); cos_data_int <= to_unsigned(54220,N);
          when 1522 =>   sin_data_int <= to_unsigned(11831,N); cos_data_int <= to_unsigned(54202,N);
          when 1523 =>   sin_data_int <= to_unsigned(11813,N); cos_data_int <= to_unsigned(54184,N);
          when 1524 =>   sin_data_int <= to_unsigned(11796,N); cos_data_int <= to_unsigned(54165,N);
          when 1525 =>   sin_data_int <= to_unsigned(11779,N); cos_data_int <= to_unsigned(54147,N);
          when 1526 =>   sin_data_int <= to_unsigned(11761,N); cos_data_int <= to_unsigned(54129,N);
          when 1527 =>   sin_data_int <= to_unsigned(11744,N); cos_data_int <= to_unsigned(54111,N);
          when 1528 =>   sin_data_int <= to_unsigned(11726,N); cos_data_int <= to_unsigned(54093,N);
          when 1529 =>   sin_data_int <= to_unsigned(11708,N); cos_data_int <= to_unsigned(54075,N);
          when 1530 =>   sin_data_int <= to_unsigned(11691,N); cos_data_int <= to_unsigned(54057,N);
          when 1531 =>   sin_data_int <= to_unsigned(11673,N); cos_data_int <= to_unsigned(54039,N);
          when 1532 =>   sin_data_int <= to_unsigned(11656,N); cos_data_int <= to_unsigned(54022,N);
          when 1533 =>   sin_data_int <= to_unsigned(11638,N); cos_data_int <= to_unsigned(54004,N);
          when 1534 =>   sin_data_int <= to_unsigned(11620,N); cos_data_int <= to_unsigned(53986,N);
          when 1535 =>   sin_data_int <= to_unsigned(11602,N); cos_data_int <= to_unsigned(53968,N);
          when 1536 =>   sin_data_int <= to_unsigned(11585,N); cos_data_int <= to_unsigned(53950,N);
          when 1537 =>   sin_data_int <= to_unsigned(11567,N); cos_data_int <= to_unsigned(53933,N);
          when 1538 =>   sin_data_int <= to_unsigned(11549,N); cos_data_int <= to_unsigned(53915,N);
          when 1539 =>   sin_data_int <= to_unsigned(11531,N); cos_data_int <= to_unsigned(53897,N);
          when 1540 =>   sin_data_int <= to_unsigned(11513,N); cos_data_int <= to_unsigned(53879,N);
          when 1541 =>   sin_data_int <= to_unsigned(11496,N); cos_data_int <= to_unsigned(53862,N);
          when 1542 =>   sin_data_int <= to_unsigned(11478,N); cos_data_int <= to_unsigned(53844,N);
          when 1543 =>   sin_data_int <= to_unsigned(11460,N); cos_data_int <= to_unsigned(53827,N);
          when 1544 =>   sin_data_int <= to_unsigned(11442,N); cos_data_int <= to_unsigned(53809,N);
          when 1545 =>   sin_data_int <= to_unsigned(11424,N); cos_data_int <= to_unsigned(53791,N);
          when 1546 =>   sin_data_int <= to_unsigned(11406,N); cos_data_int <= to_unsigned(53774,N);
          when 1547 =>   sin_data_int <= to_unsigned(11388,N); cos_data_int <= to_unsigned(53756,N);
          when 1548 =>   sin_data_int <= to_unsigned(11370,N); cos_data_int <= to_unsigned(53739,N);
          when 1549 =>   sin_data_int <= to_unsigned(11351,N); cos_data_int <= to_unsigned(53722,N);
          when 1550 =>   sin_data_int <= to_unsigned(11333,N); cos_data_int <= to_unsigned(53704,N);
          when 1551 =>   sin_data_int <= to_unsigned(11315,N); cos_data_int <= to_unsigned(53687,N);
          when 1552 =>   sin_data_int <= to_unsigned(11297,N); cos_data_int <= to_unsigned(53669,N);
          when 1553 =>   sin_data_int <= to_unsigned(11279,N); cos_data_int <= to_unsigned(53652,N);
          when 1554 =>   sin_data_int <= to_unsigned(11260,N); cos_data_int <= to_unsigned(53635,N);
          when 1555 =>   sin_data_int <= to_unsigned(11242,N); cos_data_int <= to_unsigned(53618,N);
          when 1556 =>   sin_data_int <= to_unsigned(11224,N); cos_data_int <= to_unsigned(53600,N);
          when 1557 =>   sin_data_int <= to_unsigned(11206,N); cos_data_int <= to_unsigned(53583,N);
          when 1558 =>   sin_data_int <= to_unsigned(11187,N); cos_data_int <= to_unsigned(53566,N);
          when 1559 =>   sin_data_int <= to_unsigned(11169,N); cos_data_int <= to_unsigned(53549,N);
          when 1560 =>   sin_data_int <= to_unsigned(11150,N); cos_data_int <= to_unsigned(53532,N);
          when 1561 =>   sin_data_int <= to_unsigned(11132,N); cos_data_int <= to_unsigned(53515,N);
          when 1562 =>   sin_data_int <= to_unsigned(11114,N); cos_data_int <= to_unsigned(53498,N);
          when 1563 =>   sin_data_int <= to_unsigned(11095,N); cos_data_int <= to_unsigned(53481,N);
          when 1564 =>   sin_data_int <= to_unsigned(11077,N); cos_data_int <= to_unsigned(53463,N);
          when 1565 =>   sin_data_int <= to_unsigned(11058,N); cos_data_int <= to_unsigned(53447,N);
          when 1566 =>   sin_data_int <= to_unsigned(11040,N); cos_data_int <= to_unsigned(53430,N);
          when 1567 =>   sin_data_int <= to_unsigned(11021,N); cos_data_int <= to_unsigned(53413,N);
          when 1568 =>   sin_data_int <= to_unsigned(11002,N); cos_data_int <= to_unsigned(53396,N);
          when 1569 =>   sin_data_int <= to_unsigned(10984,N); cos_data_int <= to_unsigned(53379,N);
          when 1570 =>   sin_data_int <= to_unsigned(10965,N); cos_data_int <= to_unsigned(53362,N);
          when 1571 =>   sin_data_int <= to_unsigned(10946,N); cos_data_int <= to_unsigned(53345,N);
          when 1572 =>   sin_data_int <= to_unsigned(10928,N); cos_data_int <= to_unsigned(53328,N);
          when 1573 =>   sin_data_int <= to_unsigned(10909,N); cos_data_int <= to_unsigned(53312,N);
          when 1574 =>   sin_data_int <= to_unsigned(10890,N); cos_data_int <= to_unsigned(53295,N);
          when 1575 =>   sin_data_int <= to_unsigned(10871,N); cos_data_int <= to_unsigned(53278,N);
          when 1576 =>   sin_data_int <= to_unsigned(10853,N); cos_data_int <= to_unsigned(53262,N);
          when 1577 =>   sin_data_int <= to_unsigned(10834,N); cos_data_int <= to_unsigned(53245,N);
          when 1578 =>   sin_data_int <= to_unsigned(10815,N); cos_data_int <= to_unsigned(53228,N);
          when 1579 =>   sin_data_int <= to_unsigned(10796,N); cos_data_int <= to_unsigned(53212,N);
          when 1580 =>   sin_data_int <= to_unsigned(10777,N); cos_data_int <= to_unsigned(53195,N);
          when 1581 =>   sin_data_int <= to_unsigned(10758,N); cos_data_int <= to_unsigned(53179,N);
          when 1582 =>   sin_data_int <= to_unsigned(10739,N); cos_data_int <= to_unsigned(53162,N);
          when 1583 =>   sin_data_int <= to_unsigned(10720,N); cos_data_int <= to_unsigned(53146,N);
          when 1584 =>   sin_data_int <= to_unsigned(10701,N); cos_data_int <= to_unsigned(53129,N);
          when 1585 =>   sin_data_int <= to_unsigned(10682,N); cos_data_int <= to_unsigned(53113,N);
          when 1586 =>   sin_data_int <= to_unsigned(10663,N); cos_data_int <= to_unsigned(53097,N);
          when 1587 =>   sin_data_int <= to_unsigned(10644,N); cos_data_int <= to_unsigned(53080,N);
          when 1588 =>   sin_data_int <= to_unsigned(10625,N); cos_data_int <= to_unsigned(53064,N);
          when 1589 =>   sin_data_int <= to_unsigned(10606,N); cos_data_int <= to_unsigned(53048,N);
          when 1590 =>   sin_data_int <= to_unsigned(10586,N); cos_data_int <= to_unsigned(53031,N);
          when 1591 =>   sin_data_int <= to_unsigned(10567,N); cos_data_int <= to_unsigned(53015,N);
          when 1592 =>   sin_data_int <= to_unsigned(10548,N); cos_data_int <= to_unsigned(52999,N);
          when 1593 =>   sin_data_int <= to_unsigned(10529,N); cos_data_int <= to_unsigned(52983,N);
          when 1594 =>   sin_data_int <= to_unsigned(10510,N); cos_data_int <= to_unsigned(52967,N);
          when 1595 =>   sin_data_int <= to_unsigned(10490,N); cos_data_int <= to_unsigned(52951,N);
          when 1596 =>   sin_data_int <= to_unsigned(10471,N); cos_data_int <= to_unsigned(52935,N);
          when 1597 =>   sin_data_int <= to_unsigned(10452,N); cos_data_int <= to_unsigned(52918,N);
          when 1598 =>   sin_data_int <= to_unsigned(10432,N); cos_data_int <= to_unsigned(52902,N);
          when 1599 =>   sin_data_int <= to_unsigned(10413,N); cos_data_int <= to_unsigned(52886,N);
          when 1600 =>   sin_data_int <= to_unsigned(10393,N); cos_data_int <= to_unsigned(52870,N);
          when 1601 =>   sin_data_int <= to_unsigned(10374,N); cos_data_int <= to_unsigned(52855,N);
          when 1602 =>   sin_data_int <= to_unsigned(10354,N); cos_data_int <= to_unsigned(52839,N);
          when 1603 =>   sin_data_int <= to_unsigned(10335,N); cos_data_int <= to_unsigned(52823,N);
          when 1604 =>   sin_data_int <= to_unsigned(10315,N); cos_data_int <= to_unsigned(52807,N);
          when 1605 =>   sin_data_int <= to_unsigned(10296,N); cos_data_int <= to_unsigned(52791,N);
          when 1606 =>   sin_data_int <= to_unsigned(10276,N); cos_data_int <= to_unsigned(52775,N);
          when 1607 =>   sin_data_int <= to_unsigned(10257,N); cos_data_int <= to_unsigned(52760,N);
          when 1608 =>   sin_data_int <= to_unsigned(10237,N); cos_data_int <= to_unsigned(52744,N);
          when 1609 =>   sin_data_int <= to_unsigned(10218,N); cos_data_int <= to_unsigned(52728,N);
          when 1610 =>   sin_data_int <= to_unsigned(10198,N); cos_data_int <= to_unsigned(52713,N);
          when 1611 =>   sin_data_int <= to_unsigned(10178,N); cos_data_int <= to_unsigned(52697,N);
          when 1612 =>   sin_data_int <= to_unsigned(10159,N); cos_data_int <= to_unsigned(52681,N);
          when 1613 =>   sin_data_int <= to_unsigned(10139,N); cos_data_int <= to_unsigned(52666,N);
          when 1614 =>   sin_data_int <= to_unsigned(10119,N); cos_data_int <= to_unsigned(52650,N);
          when 1615 =>   sin_data_int <= to_unsigned(10099,N); cos_data_int <= to_unsigned(52635,N);
          when 1616 =>   sin_data_int <= to_unsigned(10079,N); cos_data_int <= to_unsigned(52619,N);
          when 1617 =>   sin_data_int <= to_unsigned(10060,N); cos_data_int <= to_unsigned(52604,N);
          when 1618 =>   sin_data_int <= to_unsigned(10040,N); cos_data_int <= to_unsigned(52588,N);
          when 1619 =>   sin_data_int <= to_unsigned(10020,N); cos_data_int <= to_unsigned(52573,N);
          when 1620 =>   sin_data_int <= to_unsigned(10000,N); cos_data_int <= to_unsigned(52558,N);
          when 1621 =>   sin_data_int <= to_unsigned(9980,N); cos_data_int <= to_unsigned(52542,N);
          when 1622 =>   sin_data_int <= to_unsigned(9960,N); cos_data_int <= to_unsigned(52527,N);
          when 1623 =>   sin_data_int <= to_unsigned(9940,N); cos_data_int <= to_unsigned(52512,N);
          when 1624 =>   sin_data_int <= to_unsigned(9920,N); cos_data_int <= to_unsigned(52497,N);
          when 1625 =>   sin_data_int <= to_unsigned(9900,N); cos_data_int <= to_unsigned(52481,N);
          when 1626 =>   sin_data_int <= to_unsigned(9880,N); cos_data_int <= to_unsigned(52466,N);
          when 1627 =>   sin_data_int <= to_unsigned(9860,N); cos_data_int <= to_unsigned(52451,N);
          when 1628 =>   sin_data_int <= to_unsigned(9840,N); cos_data_int <= to_unsigned(52436,N);
          when 1629 =>   sin_data_int <= to_unsigned(9820,N); cos_data_int <= to_unsigned(52421,N);
          when 1630 =>   sin_data_int <= to_unsigned(9800,N); cos_data_int <= to_unsigned(52406,N);
          when 1631 =>   sin_data_int <= to_unsigned(9780,N); cos_data_int <= to_unsigned(52391,N);
          when 1632 =>   sin_data_int <= to_unsigned(9759,N); cos_data_int <= to_unsigned(52376,N);
          when 1633 =>   sin_data_int <= to_unsigned(9739,N); cos_data_int <= to_unsigned(52361,N);
          when 1634 =>   sin_data_int <= to_unsigned(9719,N); cos_data_int <= to_unsigned(52346,N);
          when 1635 =>   sin_data_int <= to_unsigned(9699,N); cos_data_int <= to_unsigned(52331,N);
          when 1636 =>   sin_data_int <= to_unsigned(9679,N); cos_data_int <= to_unsigned(52316,N);
          when 1637 =>   sin_data_int <= to_unsigned(9658,N); cos_data_int <= to_unsigned(52301,N);
          when 1638 =>   sin_data_int <= to_unsigned(9638,N); cos_data_int <= to_unsigned(52286,N);
          when 1639 =>   sin_data_int <= to_unsigned(9618,N); cos_data_int <= to_unsigned(52272,N);
          when 1640 =>   sin_data_int <= to_unsigned(9597,N); cos_data_int <= to_unsigned(52257,N);
          when 1641 =>   sin_data_int <= to_unsigned(9577,N); cos_data_int <= to_unsigned(52242,N);
          when 1642 =>   sin_data_int <= to_unsigned(9556,N); cos_data_int <= to_unsigned(52228,N);
          when 1643 =>   sin_data_int <= to_unsigned(9536,N); cos_data_int <= to_unsigned(52213,N);
          when 1644 =>   sin_data_int <= to_unsigned(9516,N); cos_data_int <= to_unsigned(52198,N);
          when 1645 =>   sin_data_int <= to_unsigned(9495,N); cos_data_int <= to_unsigned(52184,N);
          when 1646 =>   sin_data_int <= to_unsigned(9475,N); cos_data_int <= to_unsigned(52169,N);
          when 1647 =>   sin_data_int <= to_unsigned(9454,N); cos_data_int <= to_unsigned(52155,N);
          when 1648 =>   sin_data_int <= to_unsigned(9434,N); cos_data_int <= to_unsigned(52140,N);
          when 1649 =>   sin_data_int <= to_unsigned(9413,N); cos_data_int <= to_unsigned(52126,N);
          when 1650 =>   sin_data_int <= to_unsigned(9392,N); cos_data_int <= to_unsigned(52111,N);
          when 1651 =>   sin_data_int <= to_unsigned(9372,N); cos_data_int <= to_unsigned(52097,N);
          when 1652 =>   sin_data_int <= to_unsigned(9351,N); cos_data_int <= to_unsigned(52083,N);
          when 1653 =>   sin_data_int <= to_unsigned(9331,N); cos_data_int <= to_unsigned(52068,N);
          when 1654 =>   sin_data_int <= to_unsigned(9310,N); cos_data_int <= to_unsigned(52054,N);
          when 1655 =>   sin_data_int <= to_unsigned(9289,N); cos_data_int <= to_unsigned(52040,N);
          when 1656 =>   sin_data_int <= to_unsigned(9268,N); cos_data_int <= to_unsigned(52025,N);
          when 1657 =>   sin_data_int <= to_unsigned(9248,N); cos_data_int <= to_unsigned(52011,N);
          when 1658 =>   sin_data_int <= to_unsigned(9227,N); cos_data_int <= to_unsigned(51997,N);
          when 1659 =>   sin_data_int <= to_unsigned(9206,N); cos_data_int <= to_unsigned(51983,N);
          when 1660 =>   sin_data_int <= to_unsigned(9185,N); cos_data_int <= to_unsigned(51969,N);
          when 1661 =>   sin_data_int <= to_unsigned(9165,N); cos_data_int <= to_unsigned(51955,N);
          when 1662 =>   sin_data_int <= to_unsigned(9144,N); cos_data_int <= to_unsigned(51941,N);
          when 1663 =>   sin_data_int <= to_unsigned(9123,N); cos_data_int <= to_unsigned(51927,N);
          when 1664 =>   sin_data_int <= to_unsigned(9102,N); cos_data_int <= to_unsigned(51913,N);
          when 1665 =>   sin_data_int <= to_unsigned(9081,N); cos_data_int <= to_unsigned(51899,N);
          when 1666 =>   sin_data_int <= to_unsigned(9060,N); cos_data_int <= to_unsigned(51885,N);
          when 1667 =>   sin_data_int <= to_unsigned(9039,N); cos_data_int <= to_unsigned(51871,N);
          when 1668 =>   sin_data_int <= to_unsigned(9018,N); cos_data_int <= to_unsigned(51857,N);
          when 1669 =>   sin_data_int <= to_unsigned(8997,N); cos_data_int <= to_unsigned(51843,N);
          when 1670 =>   sin_data_int <= to_unsigned(8976,N); cos_data_int <= to_unsigned(51830,N);
          when 1671 =>   sin_data_int <= to_unsigned(8955,N); cos_data_int <= to_unsigned(51816,N);
          when 1672 =>   sin_data_int <= to_unsigned(8934,N); cos_data_int <= to_unsigned(51802,N);
          when 1673 =>   sin_data_int <= to_unsigned(8913,N); cos_data_int <= to_unsigned(51788,N);
          when 1674 =>   sin_data_int <= to_unsigned(8892,N); cos_data_int <= to_unsigned(51775,N);
          when 1675 =>   sin_data_int <= to_unsigned(8871,N); cos_data_int <= to_unsigned(51761,N);
          when 1676 =>   sin_data_int <= to_unsigned(8850,N); cos_data_int <= to_unsigned(51747,N);
          when 1677 =>   sin_data_int <= to_unsigned(8829,N); cos_data_int <= to_unsigned(51734,N);
          when 1678 =>   sin_data_int <= to_unsigned(8807,N); cos_data_int <= to_unsigned(51720,N);
          when 1679 =>   sin_data_int <= to_unsigned(8786,N); cos_data_int <= to_unsigned(51707,N);
          when 1680 =>   sin_data_int <= to_unsigned(8765,N); cos_data_int <= to_unsigned(51693,N);
          when 1681 =>   sin_data_int <= to_unsigned(8744,N); cos_data_int <= to_unsigned(51680,N);
          when 1682 =>   sin_data_int <= to_unsigned(8722,N); cos_data_int <= to_unsigned(51667,N);
          when 1683 =>   sin_data_int <= to_unsigned(8701,N); cos_data_int <= to_unsigned(51653,N);
          when 1684 =>   sin_data_int <= to_unsigned(8680,N); cos_data_int <= to_unsigned(51640,N);
          when 1685 =>   sin_data_int <= to_unsigned(8658,N); cos_data_int <= to_unsigned(51627,N);
          when 1686 =>   sin_data_int <= to_unsigned(8637,N); cos_data_int <= to_unsigned(51613,N);
          when 1687 =>   sin_data_int <= to_unsigned(8616,N); cos_data_int <= to_unsigned(51600,N);
          when 1688 =>   sin_data_int <= to_unsigned(8594,N); cos_data_int <= to_unsigned(51587,N);
          when 1689 =>   sin_data_int <= to_unsigned(8573,N); cos_data_int <= to_unsigned(51574,N);
          when 1690 =>   sin_data_int <= to_unsigned(8552,N); cos_data_int <= to_unsigned(51561,N);
          when 1691 =>   sin_data_int <= to_unsigned(8530,N); cos_data_int <= to_unsigned(51547,N);
          when 1692 =>   sin_data_int <= to_unsigned(8509,N); cos_data_int <= to_unsigned(51534,N);
          when 1693 =>   sin_data_int <= to_unsigned(8487,N); cos_data_int <= to_unsigned(51521,N);
          when 1694 =>   sin_data_int <= to_unsigned(8466,N); cos_data_int <= to_unsigned(51508,N);
          when 1695 =>   sin_data_int <= to_unsigned(8444,N); cos_data_int <= to_unsigned(51495,N);
          when 1696 =>   sin_data_int <= to_unsigned(8423,N); cos_data_int <= to_unsigned(51482,N);
          when 1697 =>   sin_data_int <= to_unsigned(8401,N); cos_data_int <= to_unsigned(51470,N);
          when 1698 =>   sin_data_int <= to_unsigned(8379,N); cos_data_int <= to_unsigned(51457,N);
          when 1699 =>   sin_data_int <= to_unsigned(8358,N); cos_data_int <= to_unsigned(51444,N);
          when 1700 =>   sin_data_int <= to_unsigned(8336,N); cos_data_int <= to_unsigned(51431,N);
          when 1701 =>   sin_data_int <= to_unsigned(8315,N); cos_data_int <= to_unsigned(51418,N);
          when 1702 =>   sin_data_int <= to_unsigned(8293,N); cos_data_int <= to_unsigned(51406,N);
          when 1703 =>   sin_data_int <= to_unsigned(8271,N); cos_data_int <= to_unsigned(51393,N);
          when 1704 =>   sin_data_int <= to_unsigned(8249,N); cos_data_int <= to_unsigned(51380,N);
          when 1705 =>   sin_data_int <= to_unsigned(8228,N); cos_data_int <= to_unsigned(51368,N);
          when 1706 =>   sin_data_int <= to_unsigned(8206,N); cos_data_int <= to_unsigned(51355,N);
          when 1707 =>   sin_data_int <= to_unsigned(8184,N); cos_data_int <= to_unsigned(51342,N);
          when 1708 =>   sin_data_int <= to_unsigned(8162,N); cos_data_int <= to_unsigned(51330,N);
          when 1709 =>   sin_data_int <= to_unsigned(8141,N); cos_data_int <= to_unsigned(51317,N);
          when 1710 =>   sin_data_int <= to_unsigned(8119,N); cos_data_int <= to_unsigned(51305,N);
          when 1711 =>   sin_data_int <= to_unsigned(8097,N); cos_data_int <= to_unsigned(51292,N);
          when 1712 =>   sin_data_int <= to_unsigned(8075,N); cos_data_int <= to_unsigned(51280,N);
          when 1713 =>   sin_data_int <= to_unsigned(8053,N); cos_data_int <= to_unsigned(51268,N);
          when 1714 =>   sin_data_int <= to_unsigned(8031,N); cos_data_int <= to_unsigned(51255,N);
          when 1715 =>   sin_data_int <= to_unsigned(8009,N); cos_data_int <= to_unsigned(51243,N);
          when 1716 =>   sin_data_int <= to_unsigned(7988,N); cos_data_int <= to_unsigned(51231,N);
          when 1717 =>   sin_data_int <= to_unsigned(7966,N); cos_data_int <= to_unsigned(51218,N);
          when 1718 =>   sin_data_int <= to_unsigned(7944,N); cos_data_int <= to_unsigned(51206,N);
          when 1719 =>   sin_data_int <= to_unsigned(7922,N); cos_data_int <= to_unsigned(51194,N);
          when 1720 =>   sin_data_int <= to_unsigned(7900,N); cos_data_int <= to_unsigned(51182,N);
          when 1721 =>   sin_data_int <= to_unsigned(7878,N); cos_data_int <= to_unsigned(51170,N);
          when 1722 =>   sin_data_int <= to_unsigned(7856,N); cos_data_int <= to_unsigned(51158,N);
          when 1723 =>   sin_data_int <= to_unsigned(7833,N); cos_data_int <= to_unsigned(51146,N);
          when 1724 =>   sin_data_int <= to_unsigned(7811,N); cos_data_int <= to_unsigned(51134,N);
          when 1725 =>   sin_data_int <= to_unsigned(7789,N); cos_data_int <= to_unsigned(51122,N);
          when 1726 =>   sin_data_int <= to_unsigned(7767,N); cos_data_int <= to_unsigned(51110,N);
          when 1727 =>   sin_data_int <= to_unsigned(7745,N); cos_data_int <= to_unsigned(51098,N);
          when 1728 =>   sin_data_int <= to_unsigned(7723,N); cos_data_int <= to_unsigned(51086,N);
          when 1729 =>   sin_data_int <= to_unsigned(7701,N); cos_data_int <= to_unsigned(51074,N);
          when 1730 =>   sin_data_int <= to_unsigned(7678,N); cos_data_int <= to_unsigned(51062,N);
          when 1731 =>   sin_data_int <= to_unsigned(7656,N); cos_data_int <= to_unsigned(51051,N);
          when 1732 =>   sin_data_int <= to_unsigned(7634,N); cos_data_int <= to_unsigned(51039,N);
          when 1733 =>   sin_data_int <= to_unsigned(7612,N); cos_data_int <= to_unsigned(51027,N);
          when 1734 =>   sin_data_int <= to_unsigned(7590,N); cos_data_int <= to_unsigned(51016,N);
          when 1735 =>   sin_data_int <= to_unsigned(7567,N); cos_data_int <= to_unsigned(51004,N);
          when 1736 =>   sin_data_int <= to_unsigned(7545,N); cos_data_int <= to_unsigned(50992,N);
          when 1737 =>   sin_data_int <= to_unsigned(7523,N); cos_data_int <= to_unsigned(50981,N);
          when 1738 =>   sin_data_int <= to_unsigned(7500,N); cos_data_int <= to_unsigned(50969,N);
          when 1739 =>   sin_data_int <= to_unsigned(7478,N); cos_data_int <= to_unsigned(50958,N);
          when 1740 =>   sin_data_int <= to_unsigned(7456,N); cos_data_int <= to_unsigned(50946,N);
          when 1741 =>   sin_data_int <= to_unsigned(7433,N); cos_data_int <= to_unsigned(50935,N);
          when 1742 =>   sin_data_int <= to_unsigned(7411,N); cos_data_int <= to_unsigned(50924,N);
          when 1743 =>   sin_data_int <= to_unsigned(7388,N); cos_data_int <= to_unsigned(50912,N);
          when 1744 =>   sin_data_int <= to_unsigned(7366,N); cos_data_int <= to_unsigned(50901,N);
          when 1745 =>   sin_data_int <= to_unsigned(7343,N); cos_data_int <= to_unsigned(50890,N);
          when 1746 =>   sin_data_int <= to_unsigned(7321,N); cos_data_int <= to_unsigned(50878,N);
          when 1747 =>   sin_data_int <= to_unsigned(7299,N); cos_data_int <= to_unsigned(50867,N);
          when 1748 =>   sin_data_int <= to_unsigned(7276,N); cos_data_int <= to_unsigned(50856,N);
          when 1749 =>   sin_data_int <= to_unsigned(7253,N); cos_data_int <= to_unsigned(50845,N);
          when 1750 =>   sin_data_int <= to_unsigned(7231,N); cos_data_int <= to_unsigned(50834,N);
          when 1751 =>   sin_data_int <= to_unsigned(7208,N); cos_data_int <= to_unsigned(50823,N);
          when 1752 =>   sin_data_int <= to_unsigned(7186,N); cos_data_int <= to_unsigned(50812,N);
          when 1753 =>   sin_data_int <= to_unsigned(7163,N); cos_data_int <= to_unsigned(50801,N);
          when 1754 =>   sin_data_int <= to_unsigned(7141,N); cos_data_int <= to_unsigned(50790,N);
          when 1755 =>   sin_data_int <= to_unsigned(7118,N); cos_data_int <= to_unsigned(50779,N);
          when 1756 =>   sin_data_int <= to_unsigned(7095,N); cos_data_int <= to_unsigned(50768,N);
          when 1757 =>   sin_data_int <= to_unsigned(7073,N); cos_data_int <= to_unsigned(50757,N);
          when 1758 =>   sin_data_int <= to_unsigned(7050,N); cos_data_int <= to_unsigned(50746,N);
          when 1759 =>   sin_data_int <= to_unsigned(7027,N); cos_data_int <= to_unsigned(50735,N);
          when 1760 =>   sin_data_int <= to_unsigned(7005,N); cos_data_int <= to_unsigned(50725,N);
          when 1761 =>   sin_data_int <= to_unsigned(6982,N); cos_data_int <= to_unsigned(50714,N);
          when 1762 =>   sin_data_int <= to_unsigned(6959,N); cos_data_int <= to_unsigned(50703,N);
          when 1763 =>   sin_data_int <= to_unsigned(6936,N); cos_data_int <= to_unsigned(50692,N);
          when 1764 =>   sin_data_int <= to_unsigned(6914,N); cos_data_int <= to_unsigned(50682,N);
          when 1765 =>   sin_data_int <= to_unsigned(6891,N); cos_data_int <= to_unsigned(50671,N);
          when 1766 =>   sin_data_int <= to_unsigned(6868,N); cos_data_int <= to_unsigned(50661,N);
          when 1767 =>   sin_data_int <= to_unsigned(6845,N); cos_data_int <= to_unsigned(50650,N);
          when 1768 =>   sin_data_int <= to_unsigned(6822,N); cos_data_int <= to_unsigned(50640,N);
          when 1769 =>   sin_data_int <= to_unsigned(6799,N); cos_data_int <= to_unsigned(50629,N);
          when 1770 =>   sin_data_int <= to_unsigned(6777,N); cos_data_int <= to_unsigned(50619,N);
          when 1771 =>   sin_data_int <= to_unsigned(6754,N); cos_data_int <= to_unsigned(50608,N);
          when 1772 =>   sin_data_int <= to_unsigned(6731,N); cos_data_int <= to_unsigned(50598,N);
          when 1773 =>   sin_data_int <= to_unsigned(6708,N); cos_data_int <= to_unsigned(50588,N);
          when 1774 =>   sin_data_int <= to_unsigned(6685,N); cos_data_int <= to_unsigned(50578,N);
          when 1775 =>   sin_data_int <= to_unsigned(6662,N); cos_data_int <= to_unsigned(50567,N);
          when 1776 =>   sin_data_int <= to_unsigned(6639,N); cos_data_int <= to_unsigned(50557,N);
          when 1777 =>   sin_data_int <= to_unsigned(6616,N); cos_data_int <= to_unsigned(50547,N);
          when 1778 =>   sin_data_int <= to_unsigned(6593,N); cos_data_int <= to_unsigned(50537,N);
          when 1779 =>   sin_data_int <= to_unsigned(6570,N); cos_data_int <= to_unsigned(50527,N);
          when 1780 =>   sin_data_int <= to_unsigned(6547,N); cos_data_int <= to_unsigned(50517,N);
          when 1781 =>   sin_data_int <= to_unsigned(6524,N); cos_data_int <= to_unsigned(50507,N);
          when 1782 =>   sin_data_int <= to_unsigned(6501,N); cos_data_int <= to_unsigned(50497,N);
          when 1783 =>   sin_data_int <= to_unsigned(6478,N); cos_data_int <= to_unsigned(50487,N);
          when 1784 =>   sin_data_int <= to_unsigned(6455,N); cos_data_int <= to_unsigned(50477,N);
          when 1785 =>   sin_data_int <= to_unsigned(6432,N); cos_data_int <= to_unsigned(50467,N);
          when 1786 =>   sin_data_int <= to_unsigned(6408,N); cos_data_int <= to_unsigned(50457,N);
          when 1787 =>   sin_data_int <= to_unsigned(6385,N); cos_data_int <= to_unsigned(50447,N);
          when 1788 =>   sin_data_int <= to_unsigned(6362,N); cos_data_int <= to_unsigned(50437,N);
          when 1789 =>   sin_data_int <= to_unsigned(6339,N); cos_data_int <= to_unsigned(50428,N);
          when 1790 =>   sin_data_int <= to_unsigned(6316,N); cos_data_int <= to_unsigned(50418,N);
          when 1791 =>   sin_data_int <= to_unsigned(6293,N); cos_data_int <= to_unsigned(50408,N);
          when 1792 =>   sin_data_int <= to_unsigned(6269,N); cos_data_int <= to_unsigned(50399,N);
          when 1793 =>   sin_data_int <= to_unsigned(6246,N); cos_data_int <= to_unsigned(50389,N);
          when 1794 =>   sin_data_int <= to_unsigned(6223,N); cos_data_int <= to_unsigned(50379,N);
          when 1795 =>   sin_data_int <= to_unsigned(6200,N); cos_data_int <= to_unsigned(50370,N);
          when 1796 =>   sin_data_int <= to_unsigned(6176,N); cos_data_int <= to_unsigned(50360,N);
          when 1797 =>   sin_data_int <= to_unsigned(6153,N); cos_data_int <= to_unsigned(50351,N);
          when 1798 =>   sin_data_int <= to_unsigned(6130,N); cos_data_int <= to_unsigned(50342,N);
          when 1799 =>   sin_data_int <= to_unsigned(6106,N); cos_data_int <= to_unsigned(50332,N);
          when 1800 =>   sin_data_int <= to_unsigned(6083,N); cos_data_int <= to_unsigned(50323,N);
          when 1801 =>   sin_data_int <= to_unsigned(6060,N); cos_data_int <= to_unsigned(50314,N);
          when 1802 =>   sin_data_int <= to_unsigned(6036,N); cos_data_int <= to_unsigned(50304,N);
          when 1803 =>   sin_data_int <= to_unsigned(6013,N); cos_data_int <= to_unsigned(50295,N);
          when 1804 =>   sin_data_int <= to_unsigned(5990,N); cos_data_int <= to_unsigned(50286,N);
          when 1805 =>   sin_data_int <= to_unsigned(5966,N); cos_data_int <= to_unsigned(50277,N);
          when 1806 =>   sin_data_int <= to_unsigned(5943,N); cos_data_int <= to_unsigned(50268,N);
          when 1807 =>   sin_data_int <= to_unsigned(5919,N); cos_data_int <= to_unsigned(50258,N);
          when 1808 =>   sin_data_int <= to_unsigned(5896,N); cos_data_int <= to_unsigned(50249,N);
          when 1809 =>   sin_data_int <= to_unsigned(5873,N); cos_data_int <= to_unsigned(50240,N);
          when 1810 =>   sin_data_int <= to_unsigned(5849,N); cos_data_int <= to_unsigned(50231,N);
          when 1811 =>   sin_data_int <= to_unsigned(5826,N); cos_data_int <= to_unsigned(50222,N);
          when 1812 =>   sin_data_int <= to_unsigned(5802,N); cos_data_int <= to_unsigned(50213,N);
          when 1813 =>   sin_data_int <= to_unsigned(5779,N); cos_data_int <= to_unsigned(50205,N);
          when 1814 =>   sin_data_int <= to_unsigned(5755,N); cos_data_int <= to_unsigned(50196,N);
          when 1815 =>   sin_data_int <= to_unsigned(5732,N); cos_data_int <= to_unsigned(50187,N);
          when 1816 =>   sin_data_int <= to_unsigned(5708,N); cos_data_int <= to_unsigned(50178,N);
          when 1817 =>   sin_data_int <= to_unsigned(5684,N); cos_data_int <= to_unsigned(50169,N);
          when 1818 =>   sin_data_int <= to_unsigned(5661,N); cos_data_int <= to_unsigned(50161,N);
          when 1819 =>   sin_data_int <= to_unsigned(5637,N); cos_data_int <= to_unsigned(50152,N);
          when 1820 =>   sin_data_int <= to_unsigned(5614,N); cos_data_int <= to_unsigned(50143,N);
          when 1821 =>   sin_data_int <= to_unsigned(5590,N); cos_data_int <= to_unsigned(50135,N);
          when 1822 =>   sin_data_int <= to_unsigned(5566,N); cos_data_int <= to_unsigned(50126,N);
          when 1823 =>   sin_data_int <= to_unsigned(5543,N); cos_data_int <= to_unsigned(50118,N);
          when 1824 =>   sin_data_int <= to_unsigned(5519,N); cos_data_int <= to_unsigned(50109,N);
          when 1825 =>   sin_data_int <= to_unsigned(5495,N); cos_data_int <= to_unsigned(50101,N);
          when 1826 =>   sin_data_int <= to_unsigned(5472,N); cos_data_int <= to_unsigned(50092,N);
          when 1827 =>   sin_data_int <= to_unsigned(5448,N); cos_data_int <= to_unsigned(50084,N);
          when 1828 =>   sin_data_int <= to_unsigned(5424,N); cos_data_int <= to_unsigned(50076,N);
          when 1829 =>   sin_data_int <= to_unsigned(5401,N); cos_data_int <= to_unsigned(50067,N);
          when 1830 =>   sin_data_int <= to_unsigned(5377,N); cos_data_int <= to_unsigned(50059,N);
          when 1831 =>   sin_data_int <= to_unsigned(5353,N); cos_data_int <= to_unsigned(50051,N);
          when 1832 =>   sin_data_int <= to_unsigned(5329,N); cos_data_int <= to_unsigned(50043,N);
          when 1833 =>   sin_data_int <= to_unsigned(5306,N); cos_data_int <= to_unsigned(50035,N);
          when 1834 =>   sin_data_int <= to_unsigned(5282,N); cos_data_int <= to_unsigned(50026,N);
          when 1835 =>   sin_data_int <= to_unsigned(5258,N); cos_data_int <= to_unsigned(50018,N);
          when 1836 =>   sin_data_int <= to_unsigned(5234,N); cos_data_int <= to_unsigned(50010,N);
          when 1837 =>   sin_data_int <= to_unsigned(5210,N); cos_data_int <= to_unsigned(50002,N);
          when 1838 =>   sin_data_int <= to_unsigned(5187,N); cos_data_int <= to_unsigned(49994,N);
          when 1839 =>   sin_data_int <= to_unsigned(5163,N); cos_data_int <= to_unsigned(49986,N);
          when 1840 =>   sin_data_int <= to_unsigned(5139,N); cos_data_int <= to_unsigned(49978,N);
          when 1841 =>   sin_data_int <= to_unsigned(5115,N); cos_data_int <= to_unsigned(49971,N);
          when 1842 =>   sin_data_int <= to_unsigned(5091,N); cos_data_int <= to_unsigned(49963,N);
          when 1843 =>   sin_data_int <= to_unsigned(5067,N); cos_data_int <= to_unsigned(49955,N);
          when 1844 =>   sin_data_int <= to_unsigned(5043,N); cos_data_int <= to_unsigned(49947,N);
          when 1845 =>   sin_data_int <= to_unsigned(5019,N); cos_data_int <= to_unsigned(49939,N);
          when 1846 =>   sin_data_int <= to_unsigned(4995,N); cos_data_int <= to_unsigned(49932,N);
          when 1847 =>   sin_data_int <= to_unsigned(4972,N); cos_data_int <= to_unsigned(49924,N);
          when 1848 =>   sin_data_int <= to_unsigned(4948,N); cos_data_int <= to_unsigned(49917,N);
          when 1849 =>   sin_data_int <= to_unsigned(4924,N); cos_data_int <= to_unsigned(49909,N);
          when 1850 =>   sin_data_int <= to_unsigned(4900,N); cos_data_int <= to_unsigned(49901,N);
          when 1851 =>   sin_data_int <= to_unsigned(4876,N); cos_data_int <= to_unsigned(49894,N);
          when 1852 =>   sin_data_int <= to_unsigned(4852,N); cos_data_int <= to_unsigned(49886,N);
          when 1853 =>   sin_data_int <= to_unsigned(4828,N); cos_data_int <= to_unsigned(49879,N);
          when 1854 =>   sin_data_int <= to_unsigned(4804,N); cos_data_int <= to_unsigned(49872,N);
          when 1855 =>   sin_data_int <= to_unsigned(4780,N); cos_data_int <= to_unsigned(49864,N);
          when 1856 =>   sin_data_int <= to_unsigned(4756,N); cos_data_int <= to_unsigned(49857,N);
          when 1857 =>   sin_data_int <= to_unsigned(4731,N); cos_data_int <= to_unsigned(49850,N);
          when 1858 =>   sin_data_int <= to_unsigned(4707,N); cos_data_int <= to_unsigned(49842,N);
          when 1859 =>   sin_data_int <= to_unsigned(4683,N); cos_data_int <= to_unsigned(49835,N);
          when 1860 =>   sin_data_int <= to_unsigned(4659,N); cos_data_int <= to_unsigned(49828,N);
          when 1861 =>   sin_data_int <= to_unsigned(4635,N); cos_data_int <= to_unsigned(49821,N);
          when 1862 =>   sin_data_int <= to_unsigned(4611,N); cos_data_int <= to_unsigned(49814,N);
          when 1863 =>   sin_data_int <= to_unsigned(4587,N); cos_data_int <= to_unsigned(49807,N);
          when 1864 =>   sin_data_int <= to_unsigned(4563,N); cos_data_int <= to_unsigned(49800,N);
          when 1865 =>   sin_data_int <= to_unsigned(4539,N); cos_data_int <= to_unsigned(49793,N);
          when 1866 =>   sin_data_int <= to_unsigned(4514,N); cos_data_int <= to_unsigned(49786,N);
          when 1867 =>   sin_data_int <= to_unsigned(4490,N); cos_data_int <= to_unsigned(49779,N);
          when 1868 =>   sin_data_int <= to_unsigned(4466,N); cos_data_int <= to_unsigned(49772,N);
          when 1869 =>   sin_data_int <= to_unsigned(4442,N); cos_data_int <= to_unsigned(49765,N);
          when 1870 =>   sin_data_int <= to_unsigned(4418,N); cos_data_int <= to_unsigned(49758,N);
          when 1871 =>   sin_data_int <= to_unsigned(4394,N); cos_data_int <= to_unsigned(49752,N);
          when 1872 =>   sin_data_int <= to_unsigned(4369,N); cos_data_int <= to_unsigned(49745,N);
          when 1873 =>   sin_data_int <= to_unsigned(4345,N); cos_data_int <= to_unsigned(49738,N);
          when 1874 =>   sin_data_int <= to_unsigned(4321,N); cos_data_int <= to_unsigned(49732,N);
          when 1875 =>   sin_data_int <= to_unsigned(4297,N); cos_data_int <= to_unsigned(49725,N);
          when 1876 =>   sin_data_int <= to_unsigned(4272,N); cos_data_int <= to_unsigned(49718,N);
          when 1877 =>   sin_data_int <= to_unsigned(4248,N); cos_data_int <= to_unsigned(49712,N);
          when 1878 =>   sin_data_int <= to_unsigned(4224,N); cos_data_int <= to_unsigned(49705,N);
          when 1879 =>   sin_data_int <= to_unsigned(4200,N); cos_data_int <= to_unsigned(49699,N);
          when 1880 =>   sin_data_int <= to_unsigned(4175,N); cos_data_int <= to_unsigned(49693,N);
          when 1881 =>   sin_data_int <= to_unsigned(4151,N); cos_data_int <= to_unsigned(49686,N);
          when 1882 =>   sin_data_int <= to_unsigned(4127,N); cos_data_int <= to_unsigned(49680,N);
          when 1883 =>   sin_data_int <= to_unsigned(4102,N); cos_data_int <= to_unsigned(49674,N);
          when 1884 =>   sin_data_int <= to_unsigned(4078,N); cos_data_int <= to_unsigned(49667,N);
          when 1885 =>   sin_data_int <= to_unsigned(4054,N); cos_data_int <= to_unsigned(49661,N);
          when 1886 =>   sin_data_int <= to_unsigned(4029,N); cos_data_int <= to_unsigned(49655,N);
          when 1887 =>   sin_data_int <= to_unsigned(4005,N); cos_data_int <= to_unsigned(49649,N);
          when 1888 =>   sin_data_int <= to_unsigned(3980,N); cos_data_int <= to_unsigned(49643,N);
          when 1889 =>   sin_data_int <= to_unsigned(3956,N); cos_data_int <= to_unsigned(49636,N);
          when 1890 =>   sin_data_int <= to_unsigned(3932,N); cos_data_int <= to_unsigned(49630,N);
          when 1891 =>   sin_data_int <= to_unsigned(3907,N); cos_data_int <= to_unsigned(49624,N);
          when 1892 =>   sin_data_int <= to_unsigned(3883,N); cos_data_int <= to_unsigned(49618,N);
          when 1893 =>   sin_data_int <= to_unsigned(3858,N); cos_data_int <= to_unsigned(49612,N);
          when 1894 =>   sin_data_int <= to_unsigned(3834,N); cos_data_int <= to_unsigned(49607,N);
          when 1895 =>   sin_data_int <= to_unsigned(3810,N); cos_data_int <= to_unsigned(49601,N);
          when 1896 =>   sin_data_int <= to_unsigned(3785,N); cos_data_int <= to_unsigned(49595,N);
          when 1897 =>   sin_data_int <= to_unsigned(3761,N); cos_data_int <= to_unsigned(49589,N);
          when 1898 =>   sin_data_int <= to_unsigned(3736,N); cos_data_int <= to_unsigned(49583,N);
          when 1899 =>   sin_data_int <= to_unsigned(3712,N); cos_data_int <= to_unsigned(49578,N);
          when 1900 =>   sin_data_int <= to_unsigned(3687,N); cos_data_int <= to_unsigned(49572,N);
          when 1901 =>   sin_data_int <= to_unsigned(3663,N); cos_data_int <= to_unsigned(49566,N);
          when 1902 =>   sin_data_int <= to_unsigned(3638,N); cos_data_int <= to_unsigned(49561,N);
          when 1903 =>   sin_data_int <= to_unsigned(3614,N); cos_data_int <= to_unsigned(49555,N);
          when 1904 =>   sin_data_int <= to_unsigned(3589,N); cos_data_int <= to_unsigned(49550,N);
          when 1905 =>   sin_data_int <= to_unsigned(3565,N); cos_data_int <= to_unsigned(49544,N);
          when 1906 =>   sin_data_int <= to_unsigned(3540,N); cos_data_int <= to_unsigned(49539,N);
          when 1907 =>   sin_data_int <= to_unsigned(3516,N); cos_data_int <= to_unsigned(49533,N);
          when 1908 =>   sin_data_int <= to_unsigned(3491,N); cos_data_int <= to_unsigned(49528,N);
          when 1909 =>   sin_data_int <= to_unsigned(3467,N); cos_data_int <= to_unsigned(49523,N);
          when 1910 =>   sin_data_int <= to_unsigned(3442,N); cos_data_int <= to_unsigned(49517,N);
          when 1911 =>   sin_data_int <= to_unsigned(3417,N); cos_data_int <= to_unsigned(49512,N);
          when 1912 =>   sin_data_int <= to_unsigned(3393,N); cos_data_int <= to_unsigned(49507,N);
          when 1913 =>   sin_data_int <= to_unsigned(3368,N); cos_data_int <= to_unsigned(49502,N);
          when 1914 =>   sin_data_int <= to_unsigned(3344,N); cos_data_int <= to_unsigned(49496,N);
          when 1915 =>   sin_data_int <= to_unsigned(3319,N); cos_data_int <= to_unsigned(49491,N);
          when 1916 =>   sin_data_int <= to_unsigned(3294,N); cos_data_int <= to_unsigned(49486,N);
          when 1917 =>   sin_data_int <= to_unsigned(3270,N); cos_data_int <= to_unsigned(49481,N);
          when 1918 =>   sin_data_int <= to_unsigned(3245,N); cos_data_int <= to_unsigned(49476,N);
          when 1919 =>   sin_data_int <= to_unsigned(3221,N); cos_data_int <= to_unsigned(49471,N);
          when 1920 =>   sin_data_int <= to_unsigned(3196,N); cos_data_int <= to_unsigned(49466,N);
          when 1921 =>   sin_data_int <= to_unsigned(3171,N); cos_data_int <= to_unsigned(49461,N);
          when 1922 =>   sin_data_int <= to_unsigned(3147,N); cos_data_int <= to_unsigned(49457,N);
          when 1923 =>   sin_data_int <= to_unsigned(3122,N); cos_data_int <= to_unsigned(49452,N);
          when 1924 =>   sin_data_int <= to_unsigned(3097,N); cos_data_int <= to_unsigned(49447,N);
          when 1925 =>   sin_data_int <= to_unsigned(3073,N); cos_data_int <= to_unsigned(49442,N);
          when 1926 =>   sin_data_int <= to_unsigned(3048,N); cos_data_int <= to_unsigned(49438,N);
          when 1927 =>   sin_data_int <= to_unsigned(3023,N); cos_data_int <= to_unsigned(49433,N);
          when 1928 =>   sin_data_int <= to_unsigned(2998,N); cos_data_int <= to_unsigned(49428,N);
          when 1929 =>   sin_data_int <= to_unsigned(2974,N); cos_data_int <= to_unsigned(49424,N);
          when 1930 =>   sin_data_int <= to_unsigned(2949,N); cos_data_int <= to_unsigned(49419,N);
          when 1931 =>   sin_data_int <= to_unsigned(2924,N); cos_data_int <= to_unsigned(49415,N);
          when 1932 =>   sin_data_int <= to_unsigned(2900,N); cos_data_int <= to_unsigned(49410,N);
          when 1933 =>   sin_data_int <= to_unsigned(2875,N); cos_data_int <= to_unsigned(49406,N);
          when 1934 =>   sin_data_int <= to_unsigned(2850,N); cos_data_int <= to_unsigned(49401,N);
          when 1935 =>   sin_data_int <= to_unsigned(2825,N); cos_data_int <= to_unsigned(49397,N);
          when 1936 =>   sin_data_int <= to_unsigned(2801,N); cos_data_int <= to_unsigned(49393,N);
          when 1937 =>   sin_data_int <= to_unsigned(2776,N); cos_data_int <= to_unsigned(49388,N);
          when 1938 =>   sin_data_int <= to_unsigned(2751,N); cos_data_int <= to_unsigned(49384,N);
          when 1939 =>   sin_data_int <= to_unsigned(2726,N); cos_data_int <= to_unsigned(49380,N);
          when 1940 =>   sin_data_int <= to_unsigned(2701,N); cos_data_int <= to_unsigned(49376,N);
          when 1941 =>   sin_data_int <= to_unsigned(2677,N); cos_data_int <= to_unsigned(49372,N);
          when 1942 =>   sin_data_int <= to_unsigned(2652,N); cos_data_int <= to_unsigned(49368,N);
          when 1943 =>   sin_data_int <= to_unsigned(2627,N); cos_data_int <= to_unsigned(49364,N);
          when 1944 =>   sin_data_int <= to_unsigned(2602,N); cos_data_int <= to_unsigned(49360,N);
          when 1945 =>   sin_data_int <= to_unsigned(2577,N); cos_data_int <= to_unsigned(49356,N);
          when 1946 =>   sin_data_int <= to_unsigned(2553,N); cos_data_int <= to_unsigned(49352,N);
          when 1947 =>   sin_data_int <= to_unsigned(2528,N); cos_data_int <= to_unsigned(49348,N);
          when 1948 =>   sin_data_int <= to_unsigned(2503,N); cos_data_int <= to_unsigned(49344,N);
          when 1949 =>   sin_data_int <= to_unsigned(2478,N); cos_data_int <= to_unsigned(49340,N);
          when 1950 =>   sin_data_int <= to_unsigned(2453,N); cos_data_int <= to_unsigned(49336,N);
          when 1951 =>   sin_data_int <= to_unsigned(2428,N); cos_data_int <= to_unsigned(49333,N);
          when 1952 =>   sin_data_int <= to_unsigned(2404,N); cos_data_int <= to_unsigned(49329,N);
          when 1953 =>   sin_data_int <= to_unsigned(2379,N); cos_data_int <= to_unsigned(49325,N);
          when 1954 =>   sin_data_int <= to_unsigned(2354,N); cos_data_int <= to_unsigned(49322,N);
          when 1955 =>   sin_data_int <= to_unsigned(2329,N); cos_data_int <= to_unsigned(49318,N);
          when 1956 =>   sin_data_int <= to_unsigned(2304,N); cos_data_int <= to_unsigned(49314,N);
          when 1957 =>   sin_data_int <= to_unsigned(2279,N); cos_data_int <= to_unsigned(49311,N);
          when 1958 =>   sin_data_int <= to_unsigned(2254,N); cos_data_int <= to_unsigned(49307,N);
          when 1959 =>   sin_data_int <= to_unsigned(2229,N); cos_data_int <= to_unsigned(49304,N);
          when 1960 =>   sin_data_int <= to_unsigned(2204,N); cos_data_int <= to_unsigned(49301,N);
          when 1961 =>   sin_data_int <= to_unsigned(2180,N); cos_data_int <= to_unsigned(49297,N);
          when 1962 =>   sin_data_int <= to_unsigned(2155,N); cos_data_int <= to_unsigned(49294,N);
          when 1963 =>   sin_data_int <= to_unsigned(2130,N); cos_data_int <= to_unsigned(49291,N);
          when 1964 =>   sin_data_int <= to_unsigned(2105,N); cos_data_int <= to_unsigned(49287,N);
          when 1965 =>   sin_data_int <= to_unsigned(2080,N); cos_data_int <= to_unsigned(49284,N);
          when 1966 =>   sin_data_int <= to_unsigned(2055,N); cos_data_int <= to_unsigned(49281,N);
          when 1967 =>   sin_data_int <= to_unsigned(2030,N); cos_data_int <= to_unsigned(49278,N);
          when 1968 =>   sin_data_int <= to_unsigned(2005,N); cos_data_int <= to_unsigned(49275,N);
          when 1969 =>   sin_data_int <= to_unsigned(1980,N); cos_data_int <= to_unsigned(49272,N);
          when 1970 =>   sin_data_int <= to_unsigned(1955,N); cos_data_int <= to_unsigned(49269,N);
          when 1971 =>   sin_data_int <= to_unsigned(1930,N); cos_data_int <= to_unsigned(49266,N);
          when 1972 =>   sin_data_int <= to_unsigned(1905,N); cos_data_int <= to_unsigned(49263,N);
          when 1973 =>   sin_data_int <= to_unsigned(1880,N); cos_data_int <= to_unsigned(49260,N);
          when 1974 =>   sin_data_int <= to_unsigned(1855,N); cos_data_int <= to_unsigned(49257,N);
          when 1975 =>   sin_data_int <= to_unsigned(1830,N); cos_data_int <= to_unsigned(49254,N);
          when 1976 =>   sin_data_int <= to_unsigned(1805,N); cos_data_int <= to_unsigned(49251,N);
          when 1977 =>   sin_data_int <= to_unsigned(1780,N); cos_data_int <= to_unsigned(49249,N);
          when 1978 =>   sin_data_int <= to_unsigned(1755,N); cos_data_int <= to_unsigned(49246,N);
          when 1979 =>   sin_data_int <= to_unsigned(1730,N); cos_data_int <= to_unsigned(49243,N);
          when 1980 =>   sin_data_int <= to_unsigned(1705,N); cos_data_int <= to_unsigned(49241,N);
          when 1981 =>   sin_data_int <= to_unsigned(1680,N); cos_data_int <= to_unsigned(49238,N);
          when 1982 =>   sin_data_int <= to_unsigned(1655,N); cos_data_int <= to_unsigned(49235,N);
          when 1983 =>   sin_data_int <= to_unsigned(1630,N); cos_data_int <= to_unsigned(49233,N);
          when 1984 =>   sin_data_int <= to_unsigned(1605,N); cos_data_int <= to_unsigned(49230,N);
          when 1985 =>   sin_data_int <= to_unsigned(1580,N); cos_data_int <= to_unsigned(49228,N);
          when 1986 =>   sin_data_int <= to_unsigned(1555,N); cos_data_int <= to_unsigned(49226,N);
          when 1987 =>   sin_data_int <= to_unsigned(1530,N); cos_data_int <= to_unsigned(49223,N);
          when 1988 =>   sin_data_int <= to_unsigned(1505,N); cos_data_int <= to_unsigned(49221,N);
          when 1989 =>   sin_data_int <= to_unsigned(1480,N); cos_data_int <= to_unsigned(49219,N);
          when 1990 =>   sin_data_int <= to_unsigned(1455,N); cos_data_int <= to_unsigned(49216,N);
          when 1991 =>   sin_data_int <= to_unsigned(1430,N); cos_data_int <= to_unsigned(49214,N);
          when 1992 =>   sin_data_int <= to_unsigned(1405,N); cos_data_int <= to_unsigned(49212,N);
          when 1993 =>   sin_data_int <= to_unsigned(1380,N); cos_data_int <= to_unsigned(49210,N);
          when 1994 =>   sin_data_int <= to_unsigned(1355,N); cos_data_int <= to_unsigned(49208,N);
          when 1995 =>   sin_data_int <= to_unsigned(1330,N); cos_data_int <= to_unsigned(49206,N);
          when 1996 =>   sin_data_int <= to_unsigned(1305,N); cos_data_int <= to_unsigned(49204,N);
          when 1997 =>   sin_data_int <= to_unsigned(1280,N); cos_data_int <= to_unsigned(49202,N);
          when 1998 =>   sin_data_int <= to_unsigned(1255,N); cos_data_int <= to_unsigned(49200,N);
          when 1999 =>   sin_data_int <= to_unsigned(1230,N); cos_data_int <= to_unsigned(49198,N);
          when 2000 =>   sin_data_int <= to_unsigned(1205,N); cos_data_int <= to_unsigned(49196,N);
          when 2001 =>   sin_data_int <= to_unsigned(1180,N); cos_data_int <= to_unsigned(49194,N);
          when 2002 =>   sin_data_int <= to_unsigned(1155,N); cos_data_int <= to_unsigned(49192,N);
          when 2003 =>   sin_data_int <= to_unsigned(1130,N); cos_data_int <= to_unsigned(49191,N);
          when 2004 =>   sin_data_int <= to_unsigned(1105,N); cos_data_int <= to_unsigned(49189,N);
          when 2005 =>   sin_data_int <= to_unsigned(1079,N); cos_data_int <= to_unsigned(49187,N);
          when 2006 =>   sin_data_int <= to_unsigned(1054,N); cos_data_int <= to_unsigned(49185,N);
          when 2007 =>   sin_data_int <= to_unsigned(1029,N); cos_data_int <= to_unsigned(49184,N);
          when 2008 =>   sin_data_int <= to_unsigned(1004,N); cos_data_int <= to_unsigned(49182,N);
          when 2009 =>   sin_data_int <= to_unsigned(979,N); cos_data_int <= to_unsigned(49181,N);
          when 2010 =>   sin_data_int <= to_unsigned(954,N); cos_data_int <= to_unsigned(49179,N);
          when 2011 =>   sin_data_int <= to_unsigned(929,N); cos_data_int <= to_unsigned(49178,N);
          when 2012 =>   sin_data_int <= to_unsigned(904,N); cos_data_int <= to_unsigned(49176,N);
          when 2013 =>   sin_data_int <= to_unsigned(879,N); cos_data_int <= to_unsigned(49175,N);
          when 2014 =>   sin_data_int <= to_unsigned(854,N); cos_data_int <= to_unsigned(49174,N);
          when 2015 =>   sin_data_int <= to_unsigned(829,N); cos_data_int <= to_unsigned(49172,N);
          when 2016 =>   sin_data_int <= to_unsigned(803,N); cos_data_int <= to_unsigned(49171,N);
          when 2017 =>   sin_data_int <= to_unsigned(778,N); cos_data_int <= to_unsigned(49170,N);
          when 2018 =>   sin_data_int <= to_unsigned(753,N); cos_data_int <= to_unsigned(49169,N);
          when 2019 =>   sin_data_int <= to_unsigned(728,N); cos_data_int <= to_unsigned(49168,N);
          when 2020 =>   sin_data_int <= to_unsigned(703,N); cos_data_int <= to_unsigned(49167,N);
          when 2021 =>   sin_data_int <= to_unsigned(678,N); cos_data_int <= to_unsigned(49166,N);
          when 2022 =>   sin_data_int <= to_unsigned(653,N); cos_data_int <= to_unsigned(49165,N);
          when 2023 =>   sin_data_int <= to_unsigned(628,N); cos_data_int <= to_unsigned(49164,N);
          when 2024 =>   sin_data_int <= to_unsigned(603,N); cos_data_int <= to_unsigned(49163,N);
          when 2025 =>   sin_data_int <= to_unsigned(577,N); cos_data_int <= to_unsigned(49162,N);
          when 2026 =>   sin_data_int <= to_unsigned(552,N); cos_data_int <= to_unsigned(49161,N);
          when 2027 =>   sin_data_int <= to_unsigned(527,N); cos_data_int <= to_unsigned(49160,N);
          when 2028 =>   sin_data_int <= to_unsigned(502,N); cos_data_int <= to_unsigned(49159,N);
          when 2029 =>   sin_data_int <= to_unsigned(477,N); cos_data_int <= to_unsigned(49158,N);
          when 2030 =>   sin_data_int <= to_unsigned(452,N); cos_data_int <= to_unsigned(49158,N);
          when 2031 =>   sin_data_int <= to_unsigned(427,N); cos_data_int <= to_unsigned(49157,N);
          when 2032 =>   sin_data_int <= to_unsigned(402,N); cos_data_int <= to_unsigned(49156,N);
          when 2033 =>   sin_data_int <= to_unsigned(376,N); cos_data_int <= to_unsigned(49156,N);
          when 2034 =>   sin_data_int <= to_unsigned(351,N); cos_data_int <= to_unsigned(49155,N);
          when 2035 =>   sin_data_int <= to_unsigned(326,N); cos_data_int <= to_unsigned(49155,N);
          when 2036 =>   sin_data_int <= to_unsigned(301,N); cos_data_int <= to_unsigned(49154,N);
          when 2037 =>   sin_data_int <= to_unsigned(276,N); cos_data_int <= to_unsigned(49154,N);
          when 2038 =>   sin_data_int <= to_unsigned(251,N); cos_data_int <= to_unsigned(49153,N);
          when 2039 =>   sin_data_int <= to_unsigned(226,N); cos_data_int <= to_unsigned(49153,N);
          when 2040 =>   sin_data_int <= to_unsigned(201,N); cos_data_int <= to_unsigned(49153,N);
          when 2041 =>   sin_data_int <= to_unsigned(175,N); cos_data_int <= to_unsigned(49152,N);
          when 2042 =>   sin_data_int <= to_unsigned(150,N); cos_data_int <= to_unsigned(49152,N);
          when 2043 =>   sin_data_int <= to_unsigned(125,N); cos_data_int <= to_unsigned(49152,N);
          when 2044 =>   sin_data_int <= to_unsigned(100,N); cos_data_int <= to_unsigned(49152,N);
          when 2045 =>   sin_data_int <= to_unsigned(75,N); cos_data_int <= to_unsigned(49152,N);
          when 2046 =>   sin_data_int <= to_unsigned(50,N); cos_data_int <= to_unsigned(49152,N);
          when 2047 =>   sin_data_int <= to_unsigned(25,N); cos_data_int <= to_unsigned(49152,N);
          when others       => null;
        end case;
      end if;
    end if;
  end process;

end rtl;
